
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd
.param width_P=2*width_N
.param width_N=3*LAMBDA

Vdd	vdd	gnd	'SUPPLY'
VX1 a0 gnd 1.8
VX2 a1 gnd 1.8
VX3 a2 gnd 0
VX4 a3 gnd 0
VX11 b0 gnd pulse 0 1.8 0ns 100ps 100ps 15ns 30ns
VX21 b1 gnd 0
VX31 b2 gnd 1.8
VX41 b3 gnd 1.8
VX0 c0 gnd 0

* SPICE3 file created from adder.ext - technology: scmos

.option scale=90n

M1000 B3N1 B3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1001 I3 OK vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1002 AW P2 NT Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1003 S3 S3N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1004 Z0 P0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1005 B1N1 B1 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1006 P0 X0 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1007 gnd P1 U1 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1008 P0N1 P0 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1009 S1 S1N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1010 S3 S3N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1011 X3 B3 A3 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1012 AF P1 vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1013 A2N1 A2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1014 OK OJ gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1015 KC G1 V2 vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1016 6R LT gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1017 S0N C0 P0 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1018 S0 S0N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1019 A1N1 A1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1020 S1 S1N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1021 gnd KP C3 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1022 S2N C2N1 P2N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1023 gnd P2 U2 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1024 gnd A3 K4 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1025 P1 X1 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1026 LT P3 vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1027 KP P1 vdd w_1336_n848# CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1028 A1N1 A1 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1029 C0N1 C0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1030 KP P2 vdd w_1336_n848# CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1031 B0N1 B0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1032 Z0 C0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1033 gnd A2 K3 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1034 B2N1 B2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1035 X3 B3N1 A3N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1036 C0N1 C0 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1037 C1 Z0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1038 C1 Z0 K0 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1039 KP C1 UP Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1040 B2N1 B2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1041 S2 S2N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1042 I2 HQ OJ vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1043 Z0 C0 M0 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1044 X2 B2 A2 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1045 A0N1 A0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1046 C1N1 C1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1047 C2N C1 V1 vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1048 C4 C4N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1049 M3 A2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1050 M4 B3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1051 gnd A1 K2 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1052 P3 X3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1053 C4 C4N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1054 C2N C1 U1 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1055 X2 B2N1 A2N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1056 VE P1 GA Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1057 A0N1 A0 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1058 P1N1 P1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1059 I0 KK C3 w_1445_n857# CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1060 M3 B2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1061 P2 X2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1062 gnd G1 C2N Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1063 AW P3 gnd Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1064 L34 G2 U3 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1065 OJ HQ gnd Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1066 V1 P1 C2N vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1067 M3 B2 K3 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1068 M4 A3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1069 G2 M3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1070 V2 P2 KC vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1071 AFF AF vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1072 Y0 A0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1073 gnd G3 L34 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1074 B0N1 B0 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1075 P2N1 P2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1076 gnd P3 GA Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1077 gnd B0 N0 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1078 M2 B1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1079 I3 AFF C4N vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1080 C2 C2N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1081 S3N C3 P3 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1082 P2N1 P2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1083 KK KC vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1084 AF C1 LO Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1085 LT G1 vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1086 S1N C1 P1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1087 MP P1 UP Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1088 G1 M2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1089 M2 B1 K2 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1090 P3N1 P3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1091 X1 B1 A1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1092 KC G1 U2 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1093 I0 KP vdd w_1445_n857# CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1094 HQ L34 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1095 C1N1 C1 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1096 M4 B3 K4 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1097 LT G1 NT Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1098 Y0 B0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1099 X0 B0N1 A0N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1100 C2N1 C2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1101 gnd 6R OJ Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1102 vdd G1 V1 vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1103 gnd P0 M0 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1104 M2 A1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1105 gnd Y0 K0 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1106 P0 X0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1107 C4N OK gnd Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1108 P1N1 P1 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1109 vdd G2 V2 vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1110 X1 B1N1 A1N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1111 AF P2 vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1112 I2 6R vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1113 OK OJ vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1114 6R LT vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1115 C3N1 C3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1116 gnd G2 KC Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1117 P2 X2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1118 S0 S0N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1119 S1N C1N1 P1N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1120 MP P2 gnd Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1121 P1 X1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1122 LT P2 vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1123 X0 B0 A0 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1124 AF C1 vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1125 G2 M3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1126 Y0 A0 N0 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1127 C1 Y0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1128 B3N1 B3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1129 AFF AF gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1130 gnd P3 U3 Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1131 L34 G2 V3 vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1132 C3N1 C3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1133 AF P3 vdd vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1134 C3 KK gnd Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1135 A3N1 A3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1136 KP C1 vdd w_1336_n848# CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1137 C2 C2N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1138 G3 M4 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1139 S2 S2N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1140 A3N1 A3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1141 KK KC gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1142 G1 M2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1143 P3N1 P3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1144 gnd AFF C4N Gnd CMOSN w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1145 P0N1 P0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1146 S0N C0N1 P0N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1147 VE P2 LO Gnd CMOSN w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1148 HQ L34 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1149 S3N C3N1 P3N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1150 A2N1 A2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1151 G3 M4 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1152 P3 X3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1153 S2N C2 P2 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1154 V3 P3 L34 vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1155 B1N1 B1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1156 C2N1 C2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1157 vdd G3 V3 vdd CMOSP w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
C0 B2N1 vdd 0.094864f
C1 M3 K3 0.061857f
C2 X2 P2 0.058778f
C3 A2 gnd 0.197904f
C4 P1 C1 0.291462f
C5 m2_1691_n440# V3 9.6e-20
C6 m3_665_n303# C0 0.026959f
C7 gnd OJ 0.207735f
C8 P1 m3_1147_n367# 1.13e-19
C9 vdd m2_1184_n874# 0.008839f
C10 P2N1 m3_1314_n716# 3.33e-19
C11 gnd S3N 0.080082f
C12 vdd B3N1 0.094864f
C13 C3 C3N1 1.62e-19
C14 m2_1314_n768# m3_1314_n716# 4.06e-19
C15 G2 V2 0.055711f
C16 U3 m2_1691_n440# 9.6e-20
C17 B0 gnd 0.056518f
C18 A2N1 vdd 0.094864f
C19 A0 m2_453_n347# 3.1e-19
C20 m3_1002_n364# A1 1.13e-19
C21 vdd B1 0.179921f
C22 gnd C4N 0.207735f
C23 B3 M4 0.11336f
C24 C2 m3_1184_n519# 1.87e-19
C25 A2N1 m3_1054_n713# 3.33e-19
C26 S2N m3_1403_n733# 1.12e-19
C27 vdd m2_1246_n763# 0.00571f
C28 HQ L34 2.74e-19
C29 OK AFF 0.135198f
C30 vdd S0N 0.067556f
C31 M3 G2 0.058778f
C32 X2 vdd 0.067556f
C33 GA gnd 0.092785f
C34 m2_1002_n416# A1N1 2.88e-19
C35 vdd AFF 0.147207f
C36 gnd m2_1548_n304# 0.002765f
C37 vdd m2_1002_n416# 0.004941f
C38 m3_2106_n415# C4 1.87e-19
C39 KK w_1445_n857# 0.044302f
C40 vdd S3 0.094864f
C41 Z0 Y0 0.227363f
C42 X1 B1 0.001447f
C43 K0 gnd 0.061857f
C44 P3 P2 0.983916f
C45 gnd LT 0.056518f
C46 vdd C1N1 0.094864f
C47 P0 Z0 0.162736f
C48 MP gnd 0.092785f
C49 vdd m2_665_n355# 0.004941f
C50 m3_1002_n364# B1 0.007496f
C51 HQ I2 0.05668f
C52 vdd A3 0.4263f
C53 S1N C1N1 4.82e-19
C54 A1 M2 0.162736f
C55 VE P2 0.05668f
C56 A0 vdd 0.405391f
C57 HQ gnd 0.127318f
C58 gnd K4 0.061857f
C59 KK MP 3.8e-20
C60 U2 P2 0.041988f
C61 vdd m2_453_n347# 0.00571f
C62 m3_2106_n415# C4N 1.12e-19
C63 HQ AW 3.8e-20
C64 m2_1002_n416# m3_1002_n364# 4.06e-19
C65 P3 vdd 0.743551f
C66 gnd S1 0.072183f
C67 G1 LT 0.264241f
C68 vdd 6R 0.235619f
C69 m3_1683_n257# P3N1 3.33e-19
C70 C2N m3_1184_n519# 1.12e-19
C71 P2N1 m2_1314_n768# 2.88e-19
C72 vdd P2 0.731754f
C73 B2N1 m2_1054_n765# 0.001081f
C74 C3 gnd 0.187116f
C75 NT AW 0.092785f
C76 A2 B2 0.251497f
C77 vdd G3 0.163748f
C78 m3_1772_n274# S3 1.87e-19
C79 B1 M2 0.11336f
C80 C3 KK 0.112874f
C81 C2 m2_1246_n763# 7.05e-19
C82 P3 m3_1679_n487# 1.53e-19
C83 A2N1 m2_1054_n765# 2.88e-19
C84 K2 A1 0.055711f
C85 m2_1683_n309# m3_1683_n257# 4.06e-19
C86 K0 C1 0.061857f
C87 GA P1 0.055711f
C88 NT G1 0.055711f
C89 OK vdd 0.194108f
C90 vdd A1N1 0.094864f
C91 gnd C0N1 0.072183f
C92 m2_665_n355# P0N1 2.88e-19
C93 KP P2 7.27e-19
C94 I0 KK 0.05668f
C95 m3_1679_n487# G3 0.002413f
C96 vdd m3_1054_n713# 0.001731f
C97 V1 vdd 0.191129f
C98 m2_1683_n309# P3N1 2.88e-19
C99 gnd A1 0.056518f
C100 vdd S1N 0.067556f
C101 m3_1423_n254# A3 1.13e-19
C102 X3 B3N1 4.82e-19
C103 G2 P2 0.006818f
C104 M3 gnd 0.056518f
C105 C1 UP 0.055711f
C106 P1 MP 0.05668f
C107 M4 K4 0.061857f
C108 vdd m3_1679_n487# 0.003759f
C109 m2_1548_n304# m3_1683_n257# 0.007496f
C110 gnd A0N1 0.072183f
C111 K2 B1 0.055711f
C112 vdd X1 0.067556f
C113 m2_1423_n306# B3N1 0.001081f
C114 B1N1 B1 1.62e-19
C115 C4N C4 1.62e-19
C116 A3 A3N1 1.62e-19
C117 P1 UP 0.055711f
C118 V2 G1 0.041965f
C119 B2N1 gnd 0.072183f
C120 KP vdd 0.426126f
C121 m3_1002_n364# A1N1 3.33e-19
C122 m2_1147_n419# C1N1 0.001081f
C123 B0 X0 0.001447f
C124 B3 K4 0.055711f
C125 C0 Z0 0.11336f
C126 vdd m3_1002_n364# 0.001885f
C127 A0 Y0 0.11336f
C128 gnd B3N1 0.072183f
C129 C1 Z0 0.11336f
C130 vdd B0N1 0.094864f
C131 A2N1 gnd 0.072183f
C132 C2 P2 6.04e-19
C133 V2 KC 0.247428f
C134 U1 m2_1094_n512# 9.6e-20
C135 G2 vdd 0.197315f
C136 gnd B1 0.059283f
C137 m2_1002_n416# B1N1 0.001081f
C138 P0 M0 0.055711f
C139 C0N1 C0 1.62e-19
C140 vdd m3_1772_n274# 0.001729f
C141 gnd m2_1246_n763# 0.002765f
C142 A0 N0 0.055711f
C143 vdd P0N1 0.094864f
C144 gnd S0N 0.080082f
C145 C2N1 vdd 0.094864f
C146 X2 gnd 0.080082f
C147 B0 m2_496_n352# 3.61e-19
C148 gnd AFF 0.085941f
C149 G1 m2_1184_n874# 6.24e-19
C150 vdd m3_1423_n254# 0.001731f
C151 C2N U1 0.061857f
C152 vdd C3N1 0.094864f
C153 gnd S3 0.072183f
C154 P3 L34 0.041965f
C155 I3 C4N 0.123714f
C156 U1 gnd 0.061857f
C157 C2 vdd 0.138746f
C158 gnd C1N1 0.072183f
C159 vdd M2 0.232636f
C160 P3 X3 0.058778f
C161 KC m2_1184_n874# 0.018008f
C162 vdd m2_1054_n765# 0.004941f
C163 S2 m3_1403_n733# 1.87e-19
C164 gnd A3 0.056518f
C165 HQ OJ 0.112874f
C166 vdd A3N1 0.094864f
C167 G3 L34 0.055711f
C168 m2_1246_n763# m3_1314_n716# 0.007496f
C169 m2_1054_n765# m3_1054_n713# 4.06e-19
C170 A0 gnd 0.056518f
C171 S2N vdd 0.067556f
C172 vdd Y0 0.312741f
C173 gnd M0 0.061857f
C174 vdd m2_1147_n419# 0.004941f
C175 gnd m2_453_n347# 0.002765f
C176 P2 w_1336_n848# 0.09959f
C177 vdd P0 0.529229f
C178 6R I2 7.27e-19
C179 AF AFF 0.058778f
C180 B2 M3 0.11336f
C181 P3 gnd 0.183685f
C182 m3_730_n320# S0 1.87e-19
C183 gnd 6R 0.168434f
C184 vdd L34 0.06532f
C185 S0N C0 0.001447f
C186 P2 gnd 0.183685f
C187 C3 m2_1683_n309# 3.61e-19
C188 vdd m2_1094_n512# 0.016328f
C189 AW P3 0.05668f
C190 C3 S3N 0.001447f
C191 vdd X3 0.067556f
C192 P3 V3 0.056801f
C193 V1 m2_1094_n512# 9.6e-20
C194 B2N1 B2 1.62e-19
C195 AW P2 0.05668f
C196 gnd G3 0.072183f
C197 vdd B1N1 0.094864f
C198 B3N1 B3 1.62e-19
C199 U2 gnd 0.061857f
C200 vdd m2_1423_n306# 0.004941f
C201 KK P2 3.77e-21
C202 m3_1679_n487# L34 2.34e-20
C203 U3 P3 0.041965f
C204 C3 w_1445_n857# 0.009614f
C205 G3 V3 0.055711f
C206 U1 C1 0.041965f
C207 C2 C2N1 1.62e-19
C208 C2N vdd 0.06532f
C209 OK gnd 0.113518f
C210 gnd A1N1 0.072183f
C211 m2_665_n355# C0 3.61e-19
C212 C1 C1N1 1.62e-19
C213 vdd I2 0.149953f
C214 G1 P2 0.290858f
C215 C3 m2_1548_n304# 7.05e-19
C216 UP MP 0.092785f
C217 vdd gnd 2.57e-19
C218 V1 C2N 0.247428f
C219 P3 AF 7.27e-19
C220 NT LT 0.092785f
C221 I0 w_1445_n857# 0.026239f
C222 X1 B1N1 4.82e-19
C223 C0 M0 0.055711f
C224 P2 m3_1314_n716# 1.13e-19
C225 U1 P1 0.041988f
C226 A2 M3 0.162736f
C227 S2N C2N1 4.82e-19
C228 LO P2 0.055711f
C229 X2 B2 0.001447f
C230 gnd S1N 0.080082f
C231 vdd V3 0.191129f
C232 P2 AF 7.27e-19
C233 G2 L34 0.174647f
C234 m3_1423_n254# A3N1 3.33e-19
C235 P0 P0N1 1.62e-19
C236 A3 M4 0.162736f
C237 S0N S0 1.62e-19
C238 K3 gnd 0.061857f
C239 G1 U2 0.041965f
C240 vdd KK 0.096594f
C241 KC P2 0.041988f
C242 LO VE 0.092785f
C243 K0 Z0 0.055711f
C244 KP w_1336_n848# 0.103092f
C245 m2_665_n355# m3_665_n303# 4.06e-19
C246 S2N C2 0.001447f
C247 vdd P1N1 0.094864f
C248 gnd X1 0.080082f
C249 A3 B3 0.252419f
C250 KC U2 0.061857f
C251 KP gnd 0.055012f
C252 vdd G1 0.452846f
C253 C1 P2 0.290858f
C254 m3_1679_n487# V3 1.87e-20
C255 gnd m3_1002_n364# 1.5e-19
C256 m2_496_n352# m3_496_n300# 4.06e-19
C257 vdd m3_1314_n716# 0.001731f
C258 A2 A2N1 1.62e-19
C259 P3 P1 0.009065f
C260 V1 G1 0.055711f
C261 m2_496_n352# A0N1 2.88e-19
C262 vdd AF 0.764456f
C263 gnd B0N1 0.072183f
C264 U3 m3_1679_n487# 2.34e-20
C265 KC vdd 0.06532f
C266 G2 gnd 0.072183f
C267 P1 P2 1.967832f
C268 KP KK 0.154624f
C269 M4 G3 0.058778f
C270 vdd m3_2106_n415# 0.001729f
C271 m2_1423_n306# m3_1423_n254# 4.06e-19
C272 VE P1 0.05668f
C273 G2 V3 0.041965f
C274 N0 Y0 0.061857f
C275 gnd P0N1 0.072183f
C276 vdd C0 0.179921f
C277 K2 M2 0.061857f
C278 C2N1 gnd 0.072183f
C279 P3 m3_1683_n257# 1.13e-19
C280 I0 C3 0.123714f
C281 C1 vdd 0.672761f
C282 m3_1236_n384# S1 1.87e-19
C283 vdd m3_1147_n367# 0.001731f
C284 C2N C2 1.62e-19
C285 V1 C1 0.041965f
C286 U3 G2 0.041965f
C287 C1 S1N 0.001447f
C288 gnd C3N1 0.072183f
C289 m2_1423_n306# A3N1 2.88e-19
C290 vdd M4 0.232636f
C291 C4N AFF 0.177461f
C292 S3N S3 1.62e-19
C293 P2N1 P2 1.62e-19
C294 C2 gnd 0.128701f
C295 P1 vdd 0.627082f
C296 gnd M2 0.056518f
C297 P3 P3N1 1.62e-19
C298 vdd m3_665_n303# 0.001769f
C299 V1 P1 0.05682f
C300 gnd A3N1 0.072183f
C301 vdd B3 0.179921f
C302 I3 AFF 0.05668f
C303 KP C1 0.264241f
C304 S2N gnd 0.080082f
C305 G2 KC 0.055711f
C306 B2 vdd 0.179921f
C307 vdd m3_1683_n257# 0.001731f
C308 B2 m3_1054_n713# 0.007496f
C309 A0 B0 0.227967f
C310 P1 X1 0.058778f
C311 vdd S0 0.094864f
C312 gnd P0 0.153444f
C313 6R OJ 0.121267f
C314 B2 K3 0.055711f
C315 C2N m2_1094_n512# 0.018008f
C316 N0 gnd 0.061857f
C317 P1 KP 7.27e-19
C318 B0 m2_453_n347# 7.05e-19
C319 P2N1 vdd 0.094864f
C320 gnd L34 0.118374f
C321 G1 M2 0.058778f
C322 gnd m2_1094_n512# 0.002765f
C323 vdd m2_1314_n768# 0.004941f
C324 gnd X3 0.080082f
C325 vdd P3N1 0.094864f
C326 V3 L34 0.247428f
C327 S2 vdd 0.094864f
C328 K2 gnd 0.061857f
C329 m2_1147_n419# P1N1 2.88e-19
C330 gnd B1N1 0.072183f
C331 vdd C4 0.094864f
C332 vdd m2_1691_n440# 0.008839f
C333 P3 GA 0.055711f
C334 vdd X0 0.067556f
C335 OK OJ 0.058778f
C336 U3 L34 0.061857f
C337 P3 m2_1548_n304# 0.007565f
C338 A2 vdd 0.4263f
C339 C2N gnd 0.118374f
C340 m3_665_n303# P0N1 3.33e-19
C341 vdd OJ 0.053537f
C342 A3 K4 0.055711f
C343 A2 m3_1054_n713# 1.13e-19
C344 V2 m2_1184_n874# 9.6e-20
C345 G1 m2_1094_n512# 0.01263f
C346 vdd m2_1683_n309# 0.004941f
C347 VE GA 0.092785f
C348 OK C4N 0.056757f
C349 P3 LT 7.27e-19
C350 vdd S3N 0.067556f
C351 LT 6R 0.058778f
C352 B0 vdd 0.19512f
C353 A2 K3 0.055711f
C354 AW gnd 0.092785f
C355 C1 Y0 0.162736f
C356 vdd C4N 0.053819f
C357 m3_1423_n254# B3 0.007496f
C358 P2 LT 7.27e-19
C359 m3_496_n300# A0N1 3.33e-19
C360 P0 C0 0.243565f
C361 S0N C0N1 4.82e-19
C362 MP P2 0.05668f
C363 KK gnd 0.127206f
C364 C1 m2_1147_n419# 3.61e-19
C365 vdd m2_496_n352# 0.004941f
C366 HQ P3 9.58e-19
C367 HQ 6R 0.154624f
C368 OK I3 7.27e-19
C369 A1 B1 0.252419f
C370 m2_1147_n419# m3_1147_n367# 4.06e-19
C371 U3 gnd 0.061857f
C372 C2N G1 0.055711f
C373 gnd P1N1 0.072183f
C374 m3_730_n320# S0N 1.12e-19
C375 vdd I3 0.149953f
C376 X0 B0N1 4.82e-19
C377 G1 gnd 0.072183f
C378 vdd m2_1548_n304# 0.00571f
C379 C1 m2_1094_n512# 0.001329f
C380 B2 m2_1054_n765# 3.61e-19
C381 C2N1 m2_1314_n768# 0.001081f
C382 G2 m2_1691_n440# 6.24e-19
C383 Z0 M0 0.061857f
C384 m2_1094_n512# m3_1147_n367# 0.007496f
C385 P3 C3 6.04e-19
C386 NT P2 0.055711f
C387 m3_665_n303# P0 1.13e-19
C388 gnd AF 0.05563f
C389 vdd LT 0.518157f
C390 m2_665_n355# C0N1 0.001081f
C391 C2 m2_1314_n768# 3.61e-19
C392 KC gnd 0.118374f
C393 P1 m2_1094_n512# 0.089674f
C394 C1 w_1336_n848# 0.076833f
C395 KP w_1445_n857# 0.036219f
C396 B0 B0N1 1.62e-19
C397 X2 B2N1 4.82e-19
C398 C2N C1 0.174647f
C399 HQ vdd 0.140896f
C400 m3_1772_n274# S3N 1.12e-19
C401 gnd C0 0.05959f
C402 m2_496_n352# B0N1 0.001081f
C403 X3 B3 0.001447f
C404 C1 gnd 0.056518f
C405 KC KK 2.74e-19
C406 P1 w_1336_n848# 0.075639f
C407 vdd m3_1403_n733# 0.001729f
C408 C2N P1 0.041988f
C409 S2N S2 1.62e-19
C410 m2_1423_n306# B3 3.61e-19
C411 vdd S1 0.094864f
C412 gnd M4 0.056518f
C413 m2_1683_n309# C3N1 0.001081f
C414 S3N C3N1 4.82e-19
C415 P1 gnd 0.128701f
C416 A0 m3_496_n300# 1.13e-19
C417 KC G1 0.174647f
C418 V2 P2 0.05682f
C419 C3 vdd 0.043881f
C420 m2_1002_n416# B1 3.61e-19
C421 LO AF 0.092785f
C422 A0 A0N1 1.62e-19
C423 S1N S1 1.62e-19
C424 m2_453_n347# m3_496_n300# 0.007496f
C425 vdd m3_1184_n519# 0.001729f
C426 gnd m3_665_n303# 1.87e-20
C427 gnd B3 0.059283f
C428 vdd Z0 0.291414f
C429 P0 X0 0.058778f
C430 KP UP 0.092785f
C431 I0 vdd 0.123714f
C432 B2 gnd 0.059283f
C433 m2_1691_n440# L34 0.018008f
C434 m3_1147_n367# P1N1 3.33e-19
C435 vdd m3_1236_n384# 0.001729f
C436 LO C1 0.055711f
C437 gnd S0 0.072183f
C438 C1 AF 0.264241f
C439 P1 P1N1 1.62e-19
C440 B0 Y0 0.162736f
C441 vdd C0N1 0.094864f
C442 KP C3 0.121267f
C443 P2N1 gnd 0.072183f
C444 V2 vdd 0.191129f
C445 P1 G1 0.004789f
C446 m3_1236_n384# S1N 1.12e-19
C447 A1 A1N1 1.62e-19
C448 vdd m3_730_n320# 0.001729f
C449 B0 N0 0.055711f
C450 P1 AF 7.27e-19
C451 vdd A1 0.4263f
C452 gnd P3N1 0.072183f
C453 S2 gnd 0.072183f
C454 KP I0 7.27e-19
C455 M3 vdd 0.232635f
C456 gnd C4 0.072183f
C457 vdd m3_496_n300# 0.001731f
C458 P2 m2_1246_n763# 0.007565f
C459 U2 m2_1184_n874# 9.6e-20
C460 vdd A0N1 0.094864f
C461 K0 Y0 0.055711f
C462 gnd X0 0.080082f
C463 I2 OJ 0.123714f
C464 m3_1403_n733# 0 0.016037f
C465 m3_1314_n716# 0 0.084889f
C466 m3_1054_n713# 0 0.084889f
C467 m3_1184_n519# 0 0.016037f
C468 m3_2106_n415# 0 0.016037f
C469 m3_1679_n487# 0 0.120846f
C470 m3_1236_n384# 0 0.016037f
C471 m3_1147_n367# 0 0.084889f
C472 m3_1002_n364# 0 0.071033f
C473 m3_730_n320# 0 0.016037f
C474 m3_665_n303# 0 0.053257f
C475 m3_1772_n274# 0 0.016037f
C476 m3_496_n300# 0 0.084889f
C477 m3_1683_n257# 0 0.084889f
C478 m3_1423_n254# 0 0.084889f
C479 m2_1184_n874# 0 0.666347f
C480 m2_1314_n768# 0 0.787321f
C481 m2_1054_n765# 0 0.787321f
C482 m2_1246_n763# 0 2.01478f
C483 m2_1691_n440# 0 0.666347f
C484 m2_1147_n419# 0 0.787321f
C485 m2_1002_n416# 0 0.632543f
C486 m2_1683_n309# 0 0.787321f
C487 m2_1094_n512# 0 3.63858f
C488 m2_665_n355# 0 0.521987f
C489 m2_496_n352# 0 0.787321f
C490 m2_1423_n306# 0 0.787321f
C491 m2_453_n347# 0 1.7415f
C492 m2_1548_n304# 0 2.7555f
C493 gnd 0 3.29914f 
C494 P2 0 3.939939f 
C495 MP 0 0.080394f 
C496 KK 0 1.655338f 
C497 U2 0 0.079598f 
C498 UP 0 0.054318f 
C499 G1 0 1.335985f 
C500 vdd 0 55.54441f 
C501 C3 0 0.411508f 
C502 KC 0 0.556903f 
C503 K3 0 0.077618f 
C504 I0 0 0.067524f 
C505 C1 0 1.297105f 
C506 KP 0 1.12496f 
C507 V2 0 0.132907f 
C508 P1 0 2.801402f 
C509 G2 0 1.257262f 
C510 M3 0 0.488017f 
C511 B2 0 3.407897f 
C512 C2N1 0 0.143763f 
C513 B2N1 0 0.143763f 
C514 P2N1 0 0.041372f 
C515 C2 0 0.301065f 
C516 A2N1 0 0.041372f 
C517 S2 0 0.019328f 
C518 S2N 0 0.320702f 
C519 X2 0 0.316742f 
C520 A2 0 1.60881f 
C521 N0 0 0.077618f 
C522 U1 0 0.079598f 
C523 B0 0 1.061952f 
C524 K2 0 0.077618f 
C525 A0 0 1.339105f 
C526 GA 0 0.054318f 
C527 C2N 0 0.556903f 
C528 P3 0 3.506965f 
C529 K0 0 0.077618f 
C530 AW 0 0.080394f 
C531 VE 0 0.080394f 
C532 HQ 0 1.644708f 
C533 U3 0 0.079598f 
C534 OK 0 0.939642f 
C535 NT 0 0.054318f 
C536 LO 0 0.054318f 
C537 V1 0 0.132907f 
C538 M2 0 0.488017f 
C539 B1 0 3.319207f 
C540 C4 0 0.019328f 
C541 Y0 0 1.05481f 
C542 AFF 0 2.05961f 
C543 OJ 0 0.383004f 
C544 L34 0 0.556903f 
C545 C1N1 0 0.143763f 
C546 C4N 0 0.38067f 
C547 B1N1 0 0.143763f 
C548 M0 0 0.077618f 
C549 I3 0 0.067524f 
C550 I2 0 0.067524f 
C551 6R 0 0.754516f 
C552 LT 0 0.572436f 
C553 V3 0 0.132907f 
C554 G3 0 0.78977f 
C555 K4 0 0.077618f 
C556 P1N1 0 0.041372f 
C557 A1N1 0 0.041372f 
C558 S1 0 0.019328f 
C559 AF 0 1.0581f 
C560 S1N 0 0.320702f 
C561 Z0 0 1.66536f 
C562 C0 0 3.531337f 
C563 X1 0 0.316742f 
C564 C0N1 0 0.143763f 
C565 M4 0 0.488017f 
C566 B0N1 0 0.143763f 
C567 A1 0 1.60162f 
C568 B3 0 3.473987f 
C569 P0N1 0 0.041372f 
C570 A0N1 0 0.041372f 
C571 S0 0 0.019328f 
C572 C3N1 0 0.143763f 
C573 B3N1 0 0.143763f 
C574 P3N1 0 0.041372f 
C575 A3N1 0 0.041372f 
C576 S0N 0 0.320702f 
C577 X0 0 0.316742f 
C578 P0 0 1.67817f 
C579 S3 0 0.019328f 
C580 S3N 0 0.320702f 
C581 X3 0 0.316742f 
C582 A3 0 1.65179f 
C583 w_1445_n857# 0 1.43127f 
C584 w_1336_n848# 0 4.15822f 

.tran 1n 50n 0n
.measure tran tpd_rise
+ TRIG v(b0) VAL='SUPPLY/2' RISE=1
+ TARG v(s3) VAL='SUPPLY/2' FALL=1
.measure tran tpd_fall
+ TRIG v(b0) VAL='SUPPLY/2' FALL=1
+ TARG v(s3) VAL='SUPPLY/2' RISE=1
.measure tran total_prop_delay param='(tpd_rise+tpd_fall)/2'
.control

run
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))
set curplottitle= harshita_2023102073

plot v(b0)+2 v(a0) v(b1)+6 v(a1)+4 
plot v(b2)+2 v(a2) v(b3)+6 v(a3)+4 
plot v(s0)-2 v(s1) v(s2)+2 v(s3)+4 
plot v(c4)+2 v(b0)-2 v(s3)

;plot v(c)

.endc


