magic
tech scmos
timestamp 1732043112
<< nwell >>
rect 482 -293 506 -275
rect 571 -310 595 -292
rect 1606 -309 1692 -227
rect 1724 -314 1785 -252
rect 1847 -301 1916 -241
rect 1925 -301 1949 -283
rect 482 -345 506 -327
rect 587 -396 647 -362
rect 973 -384 1034 -322
rect 1791 -327 1815 -309
rect 1978 -310 2003 -253
rect 2024 -298 2048 -280
rect 2090 -310 2115 -253
rect 2130 -295 2154 -277
rect 1040 -397 1064 -379
rect 728 -453 788 -419
rect 1153 -452 1214 -390
rect 1310 -439 1379 -379
rect 1393 -439 1417 -421
rect 1220 -465 1244 -447
rect 1450 -448 1475 -391
rect 1489 -429 1513 -411
rect 1685 -413 1709 -395
rect 588 -532 648 -498
<< ntransistor >>
rect 552 -293 554 -287
rect 493 -304 495 -301
rect 582 -321 584 -318
rect 552 -334 554 -328
rect 1936 -312 1938 -309
rect 2035 -309 2037 -306
rect 2141 -306 2143 -303
rect 1645 -334 1647 -325
rect 1886 -326 1888 -317
rect 2000 -327 2002 -321
rect 1982 -334 1984 -328
rect 2112 -327 2114 -321
rect 2094 -334 2096 -328
rect 1765 -341 1767 -335
rect 1802 -338 1804 -335
rect 493 -356 495 -353
rect 1645 -354 1647 -345
rect 1886 -346 1888 -337
rect 1742 -354 1744 -348
rect 1765 -367 1767 -361
rect 1645 -382 1647 -373
rect 1886 -374 1888 -365
rect 1014 -411 1016 -405
rect 1051 -408 1053 -405
rect 616 -423 618 -417
rect 1645 -402 1647 -393
rect 991 -424 993 -418
rect 1014 -437 1016 -431
rect 616 -449 618 -443
rect 1696 -424 1698 -421
rect 1500 -440 1502 -437
rect 1404 -450 1406 -447
rect 1349 -464 1351 -455
rect 1472 -465 1474 -459
rect 1454 -472 1456 -466
rect 757 -480 759 -474
rect 1194 -479 1196 -473
rect 1231 -476 1233 -473
rect 1349 -484 1351 -475
rect 1171 -492 1173 -486
rect 757 -506 759 -500
rect 1194 -505 1196 -499
rect 1349 -512 1351 -503
rect 617 -559 619 -553
rect 617 -585 619 -579
<< ptransistor >>
rect 1678 -248 1680 -236
rect 1661 -268 1663 -256
rect 493 -287 495 -281
rect 1641 -282 1643 -270
rect 1749 -272 1751 -260
rect 1902 -260 1904 -248
rect 1882 -274 1884 -262
rect 1990 -271 1992 -259
rect 2102 -271 2104 -259
rect 582 -304 584 -298
rect 1622 -300 1624 -288
rect 1863 -292 1865 -280
rect 1741 -306 1743 -294
rect 1772 -306 1774 -294
rect 1936 -295 1938 -289
rect 1990 -303 1992 -291
rect 2035 -292 2037 -286
rect 2141 -289 2143 -283
rect 2102 -303 2104 -291
rect 493 -339 495 -333
rect 1802 -321 1804 -315
rect 998 -342 1000 -330
rect 608 -374 610 -368
rect 990 -376 992 -364
rect 1021 -376 1023 -364
rect 634 -390 636 -384
rect 1051 -391 1053 -385
rect 1178 -410 1180 -398
rect 1365 -398 1367 -386
rect 1345 -412 1347 -400
rect 1462 -409 1464 -397
rect 1696 -407 1698 -401
rect 749 -431 751 -425
rect 1326 -430 1328 -418
rect 775 -447 777 -441
rect 1170 -444 1172 -432
rect 1201 -444 1203 -432
rect 1404 -433 1406 -427
rect 1500 -423 1502 -417
rect 1462 -441 1464 -429
rect 1231 -459 1233 -453
rect 609 -510 611 -504
rect 635 -526 637 -520
<< ndiffusion >>
rect 547 -293 552 -287
rect 554 -293 560 -287
rect 492 -304 493 -301
rect 495 -304 496 -301
rect 581 -321 582 -318
rect 584 -321 585 -318
rect 548 -334 552 -328
rect 554 -334 560 -328
rect 1935 -312 1936 -309
rect 1938 -312 1939 -309
rect 2034 -309 2035 -306
rect 2037 -309 2038 -306
rect 2140 -306 2141 -303
rect 2143 -306 2144 -303
rect 1644 -334 1645 -325
rect 1647 -334 1648 -325
rect 1885 -326 1886 -317
rect 1888 -326 1889 -317
rect 1999 -327 2000 -321
rect 2002 -327 2003 -321
rect 1981 -334 1982 -328
rect 1984 -334 1985 -328
rect 2111 -327 2112 -321
rect 2114 -327 2115 -321
rect 2093 -334 2094 -328
rect 2096 -334 2097 -328
rect 1764 -341 1765 -335
rect 1767 -341 1768 -335
rect 1801 -338 1802 -335
rect 1804 -338 1805 -335
rect 492 -356 493 -353
rect 495 -356 496 -353
rect 1644 -354 1645 -345
rect 1647 -354 1648 -345
rect 1885 -346 1886 -337
rect 1888 -346 1889 -337
rect 1741 -354 1742 -348
rect 1744 -354 1745 -348
rect 1764 -367 1765 -361
rect 1767 -367 1768 -361
rect 1644 -382 1645 -373
rect 1647 -382 1648 -373
rect 1885 -374 1886 -365
rect 1888 -374 1889 -365
rect 1013 -411 1014 -405
rect 1016 -411 1017 -405
rect 1050 -408 1051 -405
rect 1053 -408 1054 -405
rect 615 -423 616 -417
rect 618 -423 619 -417
rect 1644 -402 1645 -393
rect 1647 -402 1648 -393
rect 990 -424 991 -418
rect 993 -424 994 -418
rect 1013 -437 1014 -431
rect 1016 -437 1017 -431
rect 615 -449 616 -443
rect 618 -449 619 -443
rect 1695 -424 1696 -421
rect 1698 -424 1699 -421
rect 1499 -440 1500 -437
rect 1502 -440 1503 -437
rect 1403 -450 1404 -447
rect 1406 -450 1407 -447
rect 1348 -464 1349 -455
rect 1351 -464 1352 -455
rect 1471 -465 1472 -459
rect 1474 -465 1475 -459
rect 1453 -472 1454 -466
rect 1456 -472 1457 -466
rect 756 -480 757 -474
rect 759 -480 760 -474
rect 1193 -479 1194 -473
rect 1196 -479 1197 -473
rect 1230 -476 1231 -473
rect 1233 -476 1234 -473
rect 1348 -484 1349 -475
rect 1351 -484 1352 -475
rect 1170 -492 1171 -486
rect 1173 -492 1174 -486
rect 756 -506 757 -500
rect 759 -506 760 -500
rect 1193 -505 1194 -499
rect 1196 -505 1197 -499
rect 1348 -512 1349 -503
rect 1351 -512 1352 -503
rect 616 -559 617 -553
rect 619 -559 620 -553
rect 616 -585 617 -579
rect 619 -585 620 -579
<< pdiffusion >>
rect 1677 -248 1678 -236
rect 1680 -248 1681 -236
rect 1660 -268 1661 -256
rect 1663 -268 1664 -256
rect 492 -287 493 -281
rect 495 -287 496 -281
rect 1640 -282 1641 -270
rect 1643 -282 1644 -270
rect 1748 -272 1749 -260
rect 1751 -272 1752 -260
rect 1901 -260 1902 -248
rect 1904 -260 1905 -248
rect 1881 -274 1882 -262
rect 1884 -274 1885 -262
rect 1989 -271 1990 -259
rect 1992 -271 1993 -259
rect 2101 -271 2102 -259
rect 2104 -271 2105 -259
rect 581 -304 582 -298
rect 584 -304 585 -298
rect 1621 -300 1622 -288
rect 1624 -300 1625 -288
rect 1862 -292 1863 -280
rect 1865 -292 1866 -280
rect 1740 -306 1741 -294
rect 1743 -306 1744 -294
rect 1771 -306 1772 -294
rect 1774 -306 1775 -294
rect 1935 -295 1936 -289
rect 1938 -295 1939 -289
rect 1989 -303 1990 -291
rect 1992 -303 1993 -291
rect 2034 -292 2035 -286
rect 2037 -292 2038 -286
rect 2140 -289 2141 -283
rect 2143 -289 2144 -283
rect 2101 -303 2102 -291
rect 2104 -303 2105 -291
rect 492 -339 493 -333
rect 495 -339 496 -333
rect 1801 -321 1802 -315
rect 1804 -321 1805 -315
rect 997 -342 998 -330
rect 1000 -342 1001 -330
rect 607 -374 608 -368
rect 610 -374 611 -368
rect 989 -376 990 -364
rect 992 -376 993 -364
rect 1020 -376 1021 -364
rect 1023 -376 1024 -364
rect 633 -390 634 -384
rect 636 -390 637 -384
rect 1050 -391 1051 -385
rect 1053 -391 1054 -385
rect 1177 -410 1178 -398
rect 1180 -410 1181 -398
rect 1364 -398 1365 -386
rect 1367 -398 1368 -386
rect 1344 -412 1345 -400
rect 1347 -412 1348 -400
rect 1461 -409 1462 -397
rect 1464 -409 1465 -397
rect 1695 -407 1696 -401
rect 1698 -407 1699 -401
rect 748 -431 749 -425
rect 751 -431 752 -425
rect 1325 -430 1326 -418
rect 1328 -430 1329 -418
rect 774 -447 775 -441
rect 777 -447 778 -441
rect 1169 -444 1170 -432
rect 1172 -444 1173 -432
rect 1200 -444 1201 -432
rect 1203 -444 1204 -432
rect 1403 -433 1404 -427
rect 1406 -433 1407 -427
rect 1499 -423 1500 -417
rect 1502 -423 1503 -417
rect 1461 -441 1462 -429
rect 1464 -441 1465 -429
rect 1230 -459 1231 -453
rect 1233 -459 1234 -453
rect 608 -510 609 -504
rect 611 -510 612 -504
rect 634 -526 635 -520
rect 637 -526 638 -520
<< ndcontact >>
rect 543 -293 547 -287
rect 560 -293 564 -287
rect 488 -305 492 -301
rect 496 -304 500 -300
rect 577 -322 581 -318
rect 585 -321 589 -317
rect 543 -334 548 -328
rect 560 -334 564 -328
rect 1931 -313 1935 -309
rect 1939 -312 1943 -308
rect 2030 -310 2034 -306
rect 2038 -309 2042 -305
rect 2136 -307 2140 -303
rect 2144 -306 2148 -302
rect 1640 -334 1644 -325
rect 1648 -334 1652 -325
rect 1881 -326 1885 -317
rect 1889 -326 1893 -317
rect 1995 -327 1999 -321
rect 2003 -327 2007 -321
rect 1977 -334 1981 -328
rect 1985 -334 1989 -328
rect 2107 -327 2111 -321
rect 2115 -327 2119 -321
rect 2089 -334 2093 -328
rect 2097 -334 2101 -328
rect 1760 -341 1764 -335
rect 1768 -341 1772 -335
rect 1797 -339 1801 -335
rect 1805 -338 1809 -334
rect 488 -357 492 -353
rect 496 -356 500 -352
rect 1640 -354 1644 -345
rect 1648 -354 1652 -345
rect 1881 -346 1885 -337
rect 1889 -346 1893 -337
rect 1737 -354 1741 -348
rect 1745 -354 1749 -348
rect 1760 -367 1764 -361
rect 1768 -367 1772 -361
rect 1640 -382 1644 -373
rect 1648 -382 1652 -373
rect 1881 -374 1885 -365
rect 1889 -374 1893 -365
rect 1009 -411 1013 -405
rect 1017 -411 1021 -405
rect 1046 -409 1050 -405
rect 1054 -408 1058 -404
rect 611 -423 615 -417
rect 619 -423 623 -417
rect 1640 -402 1644 -393
rect 1648 -402 1652 -393
rect 986 -424 990 -418
rect 994 -424 998 -418
rect 1009 -437 1013 -431
rect 1017 -437 1021 -431
rect 611 -449 615 -443
rect 619 -449 623 -443
rect 1691 -425 1695 -421
rect 1699 -424 1703 -420
rect 1495 -441 1499 -437
rect 1503 -440 1507 -436
rect 1399 -451 1403 -447
rect 1407 -450 1411 -446
rect 1344 -464 1348 -455
rect 1352 -464 1356 -455
rect 1467 -465 1471 -459
rect 1475 -465 1479 -459
rect 1449 -472 1453 -466
rect 1457 -472 1461 -466
rect 752 -480 756 -474
rect 760 -480 764 -474
rect 1189 -479 1193 -473
rect 1197 -479 1201 -473
rect 1226 -477 1230 -473
rect 1234 -476 1238 -472
rect 1344 -484 1348 -475
rect 1352 -484 1356 -475
rect 1166 -492 1170 -486
rect 1174 -492 1178 -486
rect 752 -506 756 -500
rect 760 -506 764 -500
rect 1189 -505 1193 -499
rect 1197 -505 1201 -499
rect 1344 -512 1348 -503
rect 1352 -512 1356 -503
rect 612 -559 616 -553
rect 620 -559 624 -553
rect 612 -585 616 -579
rect 620 -585 624 -579
<< pdcontact >>
rect 1673 -248 1677 -236
rect 1681 -248 1685 -236
rect 1656 -268 1660 -256
rect 1664 -268 1668 -256
rect 488 -287 492 -281
rect 496 -287 500 -281
rect 1636 -282 1640 -270
rect 1644 -282 1648 -270
rect 1744 -272 1748 -260
rect 1752 -272 1756 -260
rect 1897 -260 1901 -248
rect 1905 -260 1909 -248
rect 1877 -274 1881 -262
rect 1885 -274 1889 -262
rect 1985 -271 1989 -259
rect 1993 -271 1997 -259
rect 2097 -271 2101 -259
rect 2105 -271 2109 -259
rect 577 -304 581 -298
rect 585 -304 589 -298
rect 1617 -300 1621 -288
rect 1625 -300 1629 -288
rect 1858 -292 1862 -280
rect 1866 -292 1870 -280
rect 1736 -306 1740 -294
rect 1744 -306 1748 -294
rect 1767 -306 1771 -294
rect 1775 -306 1779 -294
rect 1931 -295 1935 -289
rect 1939 -295 1943 -289
rect 1985 -303 1989 -291
rect 1993 -303 1997 -291
rect 2030 -292 2034 -286
rect 2038 -292 2042 -286
rect 2136 -289 2140 -283
rect 2144 -289 2148 -283
rect 2097 -303 2101 -291
rect 2105 -303 2109 -291
rect 488 -339 492 -333
rect 496 -339 500 -333
rect 1797 -321 1801 -315
rect 1805 -321 1809 -315
rect 993 -342 997 -330
rect 1001 -342 1005 -330
rect 603 -374 607 -368
rect 611 -374 615 -368
rect 985 -376 989 -364
rect 993 -376 997 -364
rect 1016 -376 1020 -364
rect 1024 -376 1028 -364
rect 629 -390 633 -384
rect 637 -390 641 -384
rect 1046 -391 1050 -385
rect 1054 -391 1058 -385
rect 1173 -410 1177 -398
rect 1181 -410 1185 -398
rect 1360 -398 1364 -386
rect 1368 -398 1372 -386
rect 1340 -412 1344 -400
rect 1348 -412 1352 -400
rect 1457 -409 1461 -397
rect 1465 -409 1469 -397
rect 1691 -407 1695 -401
rect 1699 -407 1703 -401
rect 744 -431 748 -425
rect 752 -431 756 -425
rect 1321 -430 1325 -418
rect 1329 -430 1333 -418
rect 770 -447 774 -441
rect 778 -447 782 -441
rect 1165 -444 1169 -432
rect 1173 -444 1177 -432
rect 1196 -444 1200 -432
rect 1204 -444 1208 -432
rect 1399 -433 1403 -427
rect 1407 -433 1411 -427
rect 1495 -423 1499 -417
rect 1503 -423 1507 -417
rect 1457 -441 1461 -429
rect 1465 -441 1469 -429
rect 1226 -459 1230 -453
rect 1234 -459 1238 -453
rect 604 -510 608 -504
rect 612 -510 616 -504
rect 630 -526 634 -520
rect 638 -526 642 -520
<< polysilicon >>
rect 1678 -236 1680 -229
rect 1902 -248 1904 -241
rect 1661 -256 1663 -249
rect 1678 -251 1680 -248
rect 1641 -270 1643 -263
rect 1749 -260 1751 -253
rect 493 -281 495 -278
rect 552 -287 554 -284
rect 493 -301 495 -287
rect 1622 -288 1624 -281
rect 1661 -271 1663 -268
rect 1882 -262 1884 -255
rect 1990 -259 1992 -252
rect 2102 -259 2104 -252
rect 1749 -275 1751 -272
rect 1863 -280 1865 -273
rect 1902 -263 1904 -260
rect 1990 -274 1992 -271
rect 2102 -274 2104 -271
rect 1882 -277 1884 -274
rect 1641 -285 1643 -282
rect 552 -302 554 -293
rect 582 -298 584 -295
rect 1741 -294 1743 -287
rect 1772 -294 1774 -291
rect 2141 -283 2143 -280
rect 1936 -289 1938 -286
rect 1622 -303 1624 -300
rect 493 -307 495 -304
rect 582 -318 584 -304
rect 1863 -295 1865 -292
rect 1990 -291 1992 -284
rect 2035 -286 2037 -283
rect 1741 -309 1743 -306
rect 1772 -313 1774 -306
rect 1936 -309 1938 -295
rect 2102 -291 2104 -284
rect 1990 -306 1992 -303
rect 2035 -306 2037 -292
rect 2141 -303 2143 -289
rect 1802 -315 1804 -312
rect 582 -324 584 -321
rect 552 -328 554 -325
rect 493 -333 495 -330
rect 998 -330 1000 -323
rect 1645 -325 1647 -318
rect 1886 -317 1888 -310
rect 2102 -306 2104 -303
rect 2141 -309 2143 -306
rect 2035 -312 2037 -309
rect 1936 -315 1938 -312
rect 493 -346 495 -339
rect 552 -343 554 -334
rect 1645 -337 1647 -334
rect 1765 -335 1767 -328
rect 1802 -335 1804 -321
rect 2000 -321 2002 -318
rect 2112 -321 2114 -318
rect 1886 -329 1888 -326
rect 1982 -328 1984 -321
rect 2000 -334 2002 -327
rect 2094 -328 2096 -321
rect 2112 -334 2114 -327
rect 1886 -337 1888 -334
rect 1982 -337 1984 -334
rect 2094 -337 2096 -334
rect 1802 -341 1804 -338
rect 998 -345 1000 -342
rect 1645 -345 1647 -342
rect 1765 -344 1767 -341
rect 492 -350 495 -346
rect 493 -353 495 -350
rect 1742 -348 1744 -345
rect 1886 -353 1888 -346
rect 493 -359 495 -356
rect 990 -364 992 -357
rect 1645 -361 1647 -354
rect 1742 -361 1744 -354
rect 1765 -361 1767 -358
rect 1021 -364 1023 -361
rect 608 -368 610 -365
rect 608 -381 610 -374
rect 1645 -373 1647 -366
rect 1886 -365 1888 -358
rect 634 -384 636 -377
rect 990 -379 992 -376
rect 1021 -383 1023 -376
rect 1051 -385 1053 -382
rect 634 -393 636 -390
rect 1365 -386 1367 -379
rect 1765 -374 1767 -367
rect 1886 -377 1888 -374
rect 1645 -385 1647 -382
rect 1014 -405 1016 -398
rect 1051 -405 1053 -391
rect 1178 -398 1180 -391
rect 616 -417 618 -410
rect 1051 -411 1053 -408
rect 1345 -400 1347 -393
rect 1462 -397 1464 -390
rect 1645 -393 1647 -390
rect 1014 -414 1016 -411
rect 1178 -413 1180 -410
rect 991 -418 993 -415
rect 1326 -418 1328 -411
rect 1365 -401 1367 -398
rect 1696 -401 1698 -398
rect 1645 -409 1647 -402
rect 1462 -412 1464 -409
rect 1345 -415 1347 -412
rect 1500 -417 1502 -414
rect 616 -426 618 -423
rect 749 -425 751 -422
rect 991 -431 993 -424
rect 1014 -431 1016 -428
rect 749 -438 751 -431
rect 616 -443 618 -440
rect 775 -441 777 -434
rect 1170 -432 1172 -425
rect 1201 -432 1203 -429
rect 1404 -427 1406 -424
rect 1014 -444 1016 -437
rect 1326 -433 1328 -430
rect 1462 -429 1464 -422
rect 1696 -421 1698 -407
rect 1170 -447 1172 -444
rect 616 -456 618 -449
rect 775 -450 777 -447
rect 1201 -451 1203 -444
rect 1404 -447 1406 -433
rect 1500 -437 1502 -423
rect 1696 -427 1698 -424
rect 1462 -444 1464 -441
rect 1500 -443 1502 -440
rect 1231 -453 1233 -450
rect 1349 -455 1351 -448
rect 1404 -453 1406 -450
rect 757 -474 759 -467
rect 1194 -473 1196 -466
rect 1231 -473 1233 -459
rect 1472 -459 1474 -456
rect 1349 -467 1351 -464
rect 1454 -466 1456 -459
rect 1472 -472 1474 -465
rect 1349 -475 1351 -472
rect 1454 -475 1456 -472
rect 1231 -479 1233 -476
rect 757 -483 759 -480
rect 1194 -482 1196 -479
rect 1171 -486 1173 -483
rect 1349 -491 1351 -484
rect 757 -500 759 -497
rect 1171 -499 1173 -492
rect 1194 -499 1196 -496
rect 609 -504 611 -501
rect 1349 -503 1351 -496
rect 609 -517 611 -510
rect 757 -513 759 -506
rect 1194 -512 1196 -505
rect 635 -520 637 -513
rect 1349 -515 1351 -512
rect 635 -529 637 -526
rect 617 -553 619 -546
rect 617 -562 619 -559
rect 617 -579 619 -576
rect 617 -592 619 -585
<< polycontact >>
rect 1674 -233 1678 -229
rect 1898 -245 1902 -241
rect 1657 -253 1661 -249
rect 1637 -267 1641 -263
rect 1745 -257 1749 -253
rect 1878 -259 1882 -255
rect 1618 -285 1622 -281
rect 489 -298 493 -294
rect 1986 -256 1990 -252
rect 2098 -256 2102 -252
rect 1859 -277 1863 -273
rect 548 -302 552 -297
rect 1737 -291 1741 -287
rect 1986 -288 1990 -284
rect 578 -315 582 -311
rect 1932 -306 1936 -302
rect 1768 -313 1772 -309
rect 2098 -288 2102 -284
rect 2031 -303 2035 -299
rect 2137 -300 2141 -296
rect 1882 -314 1886 -310
rect 1641 -322 1645 -318
rect 994 -327 998 -323
rect 548 -343 552 -339
rect 1761 -332 1765 -328
rect 1798 -332 1802 -328
rect 1978 -325 1982 -321
rect 2090 -325 2094 -321
rect 1996 -334 2000 -330
rect 2108 -334 2112 -330
rect 488 -350 492 -346
rect 1882 -353 1886 -349
rect 986 -361 990 -357
rect 1641 -361 1645 -357
rect 1738 -361 1742 -357
rect 604 -381 608 -377
rect 1641 -370 1645 -366
rect 1882 -362 1886 -358
rect 630 -381 634 -377
rect 1017 -383 1021 -379
rect 1361 -383 1365 -379
rect 1761 -374 1765 -370
rect 1010 -402 1014 -398
rect 1047 -402 1051 -398
rect 1174 -395 1178 -391
rect 1341 -397 1345 -393
rect 612 -414 616 -410
rect 1458 -394 1462 -390
rect 1322 -415 1326 -411
rect 1641 -409 1645 -405
rect 987 -431 991 -427
rect 1166 -429 1170 -425
rect 745 -438 749 -434
rect 771 -438 775 -434
rect 1458 -426 1462 -422
rect 1010 -444 1014 -440
rect 1692 -418 1696 -414
rect 1400 -444 1404 -440
rect 612 -456 616 -452
rect 1197 -451 1201 -447
rect 1496 -434 1500 -430
rect 1345 -452 1349 -448
rect 753 -471 757 -467
rect 1190 -470 1194 -466
rect 1227 -470 1231 -466
rect 1450 -463 1454 -459
rect 1468 -472 1472 -468
rect 1345 -491 1349 -487
rect 1167 -499 1171 -495
rect 1345 -500 1349 -496
rect 605 -517 609 -513
rect 753 -513 757 -509
rect 1190 -512 1194 -508
rect 631 -517 635 -513
rect 613 -550 617 -546
rect 613 -592 617 -588
<< metal1 >>
rect 1576 -233 1674 -229
rect 473 -267 547 -262
rect 473 -294 477 -267
rect 482 -276 506 -272
rect 488 -281 492 -276
rect 543 -287 547 -267
rect 571 -293 595 -289
rect 453 -298 489 -294
rect 488 -308 492 -305
rect 482 -312 506 -308
rect 560 -311 564 -293
rect 577 -298 581 -293
rect 585 -310 589 -304
rect 560 -315 578 -311
rect 585 -314 623 -310
rect 482 -328 506 -324
rect 560 -328 564 -315
rect 585 -317 589 -314
rect 577 -325 581 -322
rect 488 -333 492 -328
rect 571 -329 595 -325
rect 488 -360 492 -357
rect 619 -358 623 -314
rect 482 -364 506 -360
rect 576 -362 623 -358
rect 576 -452 580 -362
rect 587 -381 604 -377
rect 587 -409 591 -381
rect 611 -398 615 -374
rect 619 -377 623 -362
rect 954 -327 994 -323
rect 619 -381 630 -377
rect 637 -398 641 -390
rect 954 -397 958 -327
rect 993 -354 997 -342
rect 993 -358 1020 -354
rect 993 -364 997 -358
rect 1016 -364 1020 -358
rect 985 -389 989 -376
rect 1024 -389 1028 -376
rect 1040 -380 1064 -376
rect 985 -393 1028 -389
rect 1046 -385 1050 -380
rect 1282 -383 1361 -379
rect 611 -402 641 -398
rect 921 -401 958 -397
rect 592 -414 612 -410
rect 619 -417 623 -402
rect 717 -419 764 -415
rect 611 -443 615 -423
rect 562 -456 612 -452
rect 577 -498 624 -494
rect 577 -588 581 -498
rect 588 -517 605 -513
rect 588 -545 592 -517
rect 612 -534 616 -510
rect 620 -513 624 -498
rect 717 -509 721 -419
rect 728 -438 745 -434
rect 728 -466 732 -438
rect 752 -455 756 -431
rect 760 -434 764 -419
rect 954 -427 958 -401
rect 986 -418 990 -393
rect 1017 -405 1021 -393
rect 1024 -398 1028 -393
rect 1134 -395 1174 -391
rect 1024 -402 1047 -398
rect 954 -431 987 -427
rect 1009 -431 1013 -411
rect 1046 -412 1050 -409
rect 1040 -416 1064 -412
rect 760 -438 771 -434
rect 778 -455 782 -447
rect 752 -459 782 -455
rect 733 -471 753 -467
rect 760 -474 764 -459
rect 1134 -465 1138 -395
rect 1173 -422 1177 -410
rect 1173 -426 1200 -422
rect 1173 -432 1177 -426
rect 1196 -432 1200 -426
rect 1165 -457 1169 -444
rect 1204 -457 1208 -444
rect 1220 -448 1244 -444
rect 1165 -461 1208 -457
rect 1226 -453 1230 -448
rect 1120 -469 1138 -465
rect 752 -500 756 -480
rect 1134 -495 1138 -469
rect 1166 -486 1170 -461
rect 1197 -473 1201 -461
rect 1204 -466 1208 -461
rect 1204 -470 1227 -466
rect 1134 -499 1167 -495
rect 1189 -499 1193 -479
rect 1226 -480 1230 -477
rect 1220 -484 1244 -480
rect 1292 -496 1296 -383
rect 1303 -397 1341 -393
rect 1303 -487 1307 -397
rect 1313 -415 1322 -411
rect 1313 -448 1317 -415
rect 1329 -440 1333 -430
rect 1348 -440 1352 -412
rect 1368 -440 1372 -398
rect 1425 -394 1458 -390
rect 1393 -422 1417 -418
rect 1399 -427 1403 -422
rect 1407 -440 1411 -433
rect 1425 -440 1429 -394
rect 1576 -405 1580 -233
rect 1588 -253 1657 -249
rect 1588 -366 1592 -253
rect 1599 -267 1637 -263
rect 1599 -357 1603 -267
rect 1609 -285 1618 -281
rect 1609 -318 1613 -285
rect 1625 -310 1629 -300
rect 1644 -310 1648 -282
rect 1664 -310 1668 -268
rect 1681 -310 1685 -248
rect 1829 -245 1898 -241
rect 1625 -314 1685 -310
rect 1705 -257 1745 -253
rect 1609 -322 1641 -318
rect 1648 -325 1652 -314
rect 1640 -345 1644 -334
rect 1599 -361 1641 -357
rect 1588 -370 1641 -366
rect 1648 -373 1652 -354
rect 1640 -393 1644 -382
rect 1437 -426 1458 -422
rect 1465 -429 1469 -409
rect 1489 -412 1513 -408
rect 1576 -409 1641 -405
rect 1495 -417 1499 -412
rect 1677 -414 1681 -314
rect 1705 -357 1709 -257
rect 1744 -284 1748 -272
rect 1744 -288 1771 -284
rect 1744 -294 1748 -288
rect 1767 -294 1771 -288
rect 1736 -319 1740 -306
rect 1775 -319 1779 -306
rect 1791 -310 1815 -306
rect 1736 -323 1779 -319
rect 1797 -315 1801 -310
rect 1737 -348 1741 -323
rect 1768 -335 1772 -323
rect 1775 -328 1779 -323
rect 1775 -332 1798 -328
rect 1705 -361 1738 -357
rect 1760 -361 1764 -341
rect 1797 -342 1801 -339
rect 1791 -346 1815 -342
rect 1829 -358 1833 -245
rect 1840 -259 1878 -255
rect 1840 -349 1844 -259
rect 1850 -277 1859 -273
rect 1850 -310 1854 -277
rect 1866 -302 1870 -292
rect 1885 -302 1889 -274
rect 1905 -302 1909 -260
rect 1953 -256 1986 -252
rect 2061 -256 2098 -252
rect 1925 -284 1949 -280
rect 1931 -289 1935 -284
rect 1939 -302 1943 -295
rect 1953 -302 1957 -256
rect 1965 -288 1986 -284
rect 1993 -291 1997 -271
rect 2024 -281 2048 -277
rect 1866 -306 1932 -302
rect 1939 -306 1957 -302
rect 1850 -314 1882 -310
rect 1889 -317 1893 -306
rect 1939 -308 1943 -306
rect 1931 -316 1935 -313
rect 1925 -320 1949 -316
rect 1881 -337 1885 -326
rect 1953 -337 1957 -306
rect 2030 -286 2034 -281
rect 2038 -299 2042 -292
rect 2061 -299 2065 -256
rect 2011 -303 2031 -299
rect 2038 -303 2065 -299
rect 1985 -311 1989 -303
rect 2011 -311 2014 -303
rect 2038 -305 2042 -303
rect 1985 -315 2014 -311
rect 2030 -313 2034 -310
rect 2061 -311 2065 -303
rect 2073 -288 2098 -284
rect 1965 -325 1978 -321
rect 1985 -328 1989 -315
rect 1995 -321 1999 -315
rect 2024 -317 2048 -313
rect 2061 -315 2068 -311
rect 2064 -320 2068 -315
rect 1996 -337 2000 -334
rect 1953 -341 2000 -337
rect 2073 -337 2078 -288
rect 2105 -291 2109 -271
rect 2130 -278 2154 -274
rect 2136 -283 2140 -278
rect 2118 -300 2137 -296
rect 2097 -311 2101 -303
rect 2118 -311 2122 -300
rect 2136 -310 2140 -307
rect 2097 -315 2122 -311
rect 2130 -314 2154 -310
rect 2097 -328 2101 -315
rect 2107 -321 2111 -315
rect 2108 -337 2112 -334
rect 2073 -341 2112 -337
rect 1840 -353 1882 -349
rect 1829 -362 1882 -358
rect 1889 -365 1893 -346
rect 1685 -396 1709 -392
rect 1691 -401 1695 -396
rect 1699 -414 1703 -407
rect 2073 -414 2078 -341
rect 1677 -418 1692 -414
rect 1699 -418 2078 -414
rect 1699 -420 1703 -418
rect 1691 -428 1695 -425
rect 1329 -444 1400 -440
rect 1407 -444 1429 -440
rect 1313 -452 1345 -448
rect 1352 -455 1356 -444
rect 1407 -446 1411 -444
rect 1399 -454 1403 -451
rect 1393 -458 1417 -454
rect 1344 -475 1348 -464
rect 1425 -475 1429 -444
rect 1480 -434 1496 -430
rect 1685 -432 1709 -428
rect 1457 -449 1461 -441
rect 1480 -449 1483 -434
rect 1495 -444 1499 -441
rect 1489 -448 1513 -444
rect 1457 -453 1483 -449
rect 1437 -463 1450 -459
rect 1457 -466 1461 -453
rect 1467 -459 1471 -453
rect 1468 -475 1472 -472
rect 1425 -479 1472 -475
rect 1303 -491 1345 -487
rect 1292 -500 1345 -496
rect 1352 -503 1356 -484
rect 717 -513 753 -509
rect 620 -517 631 -513
rect 638 -534 642 -526
rect 717 -534 720 -513
rect 612 -538 720 -534
rect 593 -550 613 -546
rect 620 -553 624 -538
rect 612 -579 616 -559
rect 563 -592 613 -588
<< m2contact >>
rect 587 -414 592 -409
rect 636 -407 641 -402
rect 728 -471 733 -466
rect 2064 -325 2069 -320
rect 588 -550 593 -545
<< metal2 >>
rect 536 -302 548 -297
rect 536 -317 540 -302
rect 474 -321 540 -317
rect 1757 -313 1768 -309
rect 474 -343 478 -321
rect 1757 -323 1761 -313
rect 1729 -327 1761 -323
rect 2069 -325 2090 -321
rect 1757 -332 1761 -327
rect 453 -346 478 -343
rect 496 -346 500 -339
rect 539 -343 548 -339
rect 539 -346 543 -343
rect 453 -347 488 -346
rect 474 -350 488 -347
rect 496 -350 543 -346
rect 570 -350 623 -346
rect 496 -352 500 -350
rect 570 -409 574 -350
rect 1006 -383 1017 -379
rect 1006 -393 1010 -383
rect 937 -397 1010 -393
rect 1006 -402 1010 -397
rect 570 -414 587 -409
rect 637 -466 641 -407
rect 1186 -451 1197 -447
rect 1186 -461 1190 -451
rect 1123 -465 1190 -461
rect 637 -471 728 -466
rect 1186 -470 1190 -465
rect 564 -550 588 -545
<< m123contact >>
rect 1960 -289 1965 -284
rect 1960 -326 1965 -321
rect 1432 -427 1437 -422
rect 1432 -464 1437 -459
<< metal3 >>
rect 496 -293 500 -287
rect 1717 -291 1737 -287
rect 496 -298 528 -293
rect 496 -300 500 -298
rect 524 -328 528 -298
rect 524 -334 543 -328
rect 937 -361 986 -357
rect 966 -440 970 -361
rect 1717 -370 1721 -291
rect 1960 -321 1965 -289
rect 2144 -296 2148 -289
rect 2144 -300 2154 -296
rect 2144 -302 2148 -300
rect 1805 -328 1809 -321
rect 1805 -332 1824 -328
rect 1805 -334 1809 -332
rect 1717 -374 1761 -370
rect 1820 -380 1824 -332
rect 1960 -380 1965 -326
rect 1820 -384 1965 -380
rect 1054 -398 1058 -391
rect 1054 -402 1064 -398
rect 1054 -404 1058 -402
rect 1120 -429 1166 -425
rect 966 -444 1010 -440
rect 1146 -508 1150 -429
rect 1432 -459 1437 -427
rect 1503 -430 1507 -423
rect 1503 -434 1514 -430
rect 1503 -436 1507 -434
rect 1234 -466 1238 -459
rect 1234 -470 1265 -466
rect 1234 -472 1238 -470
rect 1146 -512 1190 -508
rect 1261 -518 1265 -470
rect 1432 -518 1437 -464
rect 1261 -522 1437 -518
<< labels >>
rlabel nwell 502 -279 504 -277 1 vdd
rlabel pdcontact 488 -287 492 -281 1 vdd
rlabel nwell 502 -331 504 -329 1 vdd
rlabel pdcontact 488 -339 492 -333 1 vdd
rlabel nwell 591 -296 593 -294 1 vdd
rlabel pdcontact 577 -304 581 -298 1 vdd
rlabel ndcontact 577 -322 581 -318 1 gnd
rlabel ndcontact 488 -305 492 -301 1 gnd
rlabel ndcontact 488 -357 492 -353 1 gnd
rlabel polycontact 489 -298 493 -294 1 A0
rlabel ndcontact 496 -304 500 -300 1 A0N1
rlabel pdcontact 496 -287 500 -281 1 A0N1
rlabel polycontact 488 -350 492 -346 1 B0
rlabel ndcontact 496 -356 500 -352 1 B0N1
rlabel pdcontact 496 -339 500 -333 1 B0N1
rlabel polycontact 548 -343 552 -339 1 B0N1
rlabel ndcontact 543 -334 547 -329 1 A0N1
rlabel polycontact 548 -302 552 -297 1 B0
rlabel ndcontact 543 -293 547 -288 1 A0
rlabel ndcontact 560 -292 564 -288 1 X0
rlabel ndcontact 560 -333 564 -329 1 X0
rlabel polycontact 578 -315 582 -311 1 X0
rlabel pdcontact 585 -304 589 -298 1 P0
rlabel ndcontact 585 -321 589 -317 1 P0
rlabel pdcontact 629 -390 633 -384 1 vdd
rlabel pdcontact 603 -374 607 -368 1 vdd
rlabel ndcontact 619 -449 623 -443 1 gnd
rlabel pdcontact 630 -526 634 -520 1 vdd
rlabel pdcontact 604 -510 608 -504 1 vdd
rlabel ndcontact 620 -585 624 -579 1 gnd
rlabel pdcontact 770 -447 774 -441 1 vdd
rlabel pdcontact 744 -431 748 -425 1 vdd
rlabel ndcontact 760 -506 764 -500 1 gnd
rlabel m2contact 588 -550 592 -546 1 A0
rlabel polycontact 613 -550 617 -546 1 A0
rlabel polycontact 605 -517 609 -513 1 A0
rlabel polycontact 613 -592 617 -588 1 B0
rlabel polycontact 631 -517 635 -513 1 B0
rlabel pdcontact 612 -509 616 -505 1 Y0
rlabel pdcontact 638 -525 642 -521 1 Y0
rlabel ndcontact 620 -558 624 -554 1 Y0
rlabel ndcontact 612 -558 616 -554 1 N0
rlabel ndcontact 612 -584 616 -580 1 N0
rlabel polycontact 612 -456 616 -452 1 P0
rlabel polycontact 630 -381 634 -377 1 P0
rlabel m2contact 587 -414 591 -410 1 C0
rlabel polycontact 612 -414 616 -410 1 C0
rlabel polycontact 604 -381 608 -377 1 C0
rlabel pdcontact 611 -373 615 -369 1 Z0
rlabel pdcontact 637 -389 641 -385 1 Z0
rlabel ndcontact 619 -422 623 -418 1 Z0
rlabel ndcontact 611 -422 615 -418 1 M0
rlabel ndcontact 611 -448 615 -444 1 M0
rlabel m2contact 638 -406 640 -404 1 Z0
rlabel m2contact 728 -471 732 -467 1 Z0
rlabel polycontact 753 -471 757 -467 1 Z0
rlabel polycontact 745 -438 749 -434 1 Z0
rlabel polycontact 753 -513 757 -509 1 Y0
rlabel polycontact 771 -438 775 -434 1 Y0
rlabel ndcontact 752 -479 756 -475 1 K0
rlabel ndcontact 752 -505 756 -501 1 K0
rlabel pdcontact 778 -447 782 -443 1 C1
rlabel pdcontact 752 -430 756 -426 1 C1
rlabel ndcontact 760 -479 764 -475 1 C1
rlabel nwell 628 -369 632 -365 1 vdd
rlabel nwell 772 -428 776 -424 1 vdd
rlabel nwell 637 -508 641 -504 1 vdd
rlabel pdcontact 1001 -342 1005 -330 1 vdd
rlabel ndcontact 1017 -437 1021 -431 1 gnd
rlabel ndcontact 994 -424 998 -418 1 gnd
rlabel ndcontact 1046 -409 1050 -405 1 gnd
rlabel pdcontact 1046 -391 1050 -385 1 vdd
rlabel nwell 1060 -383 1062 -381 1 vdd
rlabel pdcontact 1054 -391 1058 -385 1 C2
rlabel ndcontact 1054 -408 1058 -404 1 C2
rlabel polycontact 1047 -402 1051 -398 1 C2N
rlabel ndcontact 1017 -411 1021 -405 1 C2N
rlabel pdcontact 1024 -373 1028 -367 1 C2N
rlabel pdcontact 985 -373 989 -367 1 C2N
rlabel ndcontact 986 -424 990 -418 1 C2N
rlabel polycontact 987 -431 991 -427 1 G1
rlabel polycontact 994 -327 998 -323 1 G1
rlabel polycontact 1017 -383 1021 -379 1 C1
rlabel polycontact 1010 -402 1014 -398 1 C1
rlabel polycontact 986 -361 990 -357 1 P1
rlabel polycontact 1010 -444 1014 -440 1 P1
rlabel ndcontact 1009 -410 1013 -406 1 U1
rlabel ndcontact 1009 -436 1013 -432 1 U1
rlabel pdcontact 993 -339 997 -335 1 V1
rlabel pdcontact 993 -373 997 -369 1 V1
rlabel pdcontact 1016 -373 1020 -369 1 V1
rlabel nwell 1018 -339 1022 -335 1 vdd
rlabel pdcontact 1181 -410 1185 -398 1 vdd
rlabel ndcontact 1197 -505 1201 -499 1 gnd
rlabel ndcontact 1174 -492 1178 -486 1 gnd
rlabel ndcontact 1226 -477 1230 -473 1 gnd
rlabel pdcontact 1226 -459 1230 -453 1 vdd
rlabel nwell 1240 -451 1242 -449 1 vdd
rlabel nwell 1198 -407 1202 -403 1 vdd
rlabel polycontact 1167 -499 1171 -495 1 G2
rlabel polycontact 1174 -395 1178 -391 1 G2
rlabel polycontact 1190 -512 1194 -508 1 P2
rlabel polycontact 1166 -429 1170 -425 1 P2
rlabel polycontact 1197 -451 1201 -447 1 G1
rlabel polycontact 1190 -470 1194 -466 1 G1
rlabel pdcontact 1173 -441 1177 -437 1 V2
rlabel pdcontact 1173 -407 1177 -403 1 V2
rlabel pdcontact 1196 -441 1200 -437 1 V2
rlabel ndcontact 1189 -478 1193 -474 1 U2
rlabel ndcontact 1189 -504 1193 -500 1 U2
rlabel pdcontact 1165 -441 1169 -435 1 KC
rlabel ndcontact 1166 -492 1170 -486 1 KC
rlabel polycontact 1227 -470 1231 -466 1 KC
rlabel pdcontact 1204 -441 1208 -435 1 KC
rlabel ndcontact 1197 -479 1201 -473 1 KC
rlabel ndcontact 1234 -476 1238 -472 1 KK
rlabel pdcontact 1234 -459 1238 -453 1 KK
rlabel pdcontact 1321 -430 1325 -418 1 vdd
rlabel pdcontact 1340 -412 1344 -400 1 vdd
rlabel pdcontact 1360 -398 1364 -386 1 vdd
rlabel ndcontact 1344 -512 1348 -503 1 gnd
rlabel polycontact 1361 -383 1365 -379 1 P2
rlabel polycontact 1345 -500 1349 -496 1 P2
rlabel polycontact 1322 -415 1326 -411 1 C1
rlabel polycontact 1345 -452 1349 -448 1 C1
rlabel polycontact 1341 -397 1345 -393 1 P1
rlabel polycontact 1345 -491 1349 -487 1 P1
rlabel ndcontact 1352 -481 1356 -477 1 MP
rlabel ndcontact 1352 -509 1356 -505 1 MP
rlabel ndcontact 1344 -483 1348 -479 1 UP
rlabel ndcontact 1344 -462 1348 -458 1 UP
rlabel pdcontact 1329 -427 1333 -423 1 KP
rlabel pdcontact 1348 -407 1352 -403 1 KP
rlabel pdcontact 1368 -394 1372 -390 1 KP
rlabel ndcontact 1352 -462 1356 -458 1 KP
rlabel pdcontact 1752 -272 1756 -260 1 vdd
rlabel ndcontact 1768 -367 1772 -361 1 gnd
rlabel ndcontact 1745 -354 1749 -348 1 gnd
rlabel ndcontact 1797 -339 1801 -335 1 gnd
rlabel pdcontact 1797 -321 1801 -315 1 vdd
rlabel nwell 1811 -313 1813 -311 1 vdd
rlabel nwell 1769 -269 1773 -265 1 vdd
rlabel polycontact 1745 -257 1749 -253 1 G3
rlabel pdcontact 1744 -269 1748 -265 1 V3
rlabel pdcontact 1744 -303 1748 -299 1 V3
rlabel pdcontact 1767 -303 1771 -299 1 V3
rlabel polycontact 1737 -291 1741 -287 1 P3
rlabel polycontact 1761 -374 1765 -370 1 P3
rlabel polycontact 1768 -313 1772 -309 1 G2
rlabel polycontact 1761 -332 1765 -328 1 G2
rlabel ndcontact 1760 -340 1764 -336 1 U3
rlabel ndcontact 1760 -366 1764 -362 1 U3
rlabel ndcontact 1805 -338 1809 -334 1 HQ
rlabel pdcontact 1805 -321 1809 -315 1 HQ
rlabel nwell 1376 -382 1378 -380 1 vdd
rlabel pdcontact 1457 -409 1461 -397 1 vdd
rlabel ndcontact 1475 -465 1479 -461 1 gnd
rlabel ndcontact 1449 -471 1453 -467 1 gnd
rlabel pdcontact 1465 -437 1469 -431 1 I0
rlabel pdcontact 1465 -406 1469 -400 1 I0
rlabel m123contact 1433 -463 1435 -460 1 KK
rlabel m123contact 1433 -426 1435 -423 1 KK
rlabel polycontact 1458 -426 1462 -422 1 KK
rlabel polycontact 1450 -463 1454 -459 1 KK
rlabel nwell 1472 -395 1474 -393 1 vdd
rlabel ndcontact 1495 -441 1499 -437 1 gnd
rlabel pdcontact 1495 -423 1499 -417 1 vdd
rlabel nwell 1509 -415 1511 -413 1 vdd
rlabel ndcontact 1457 -472 1461 -466 1 C3N
rlabel ndcontact 1467 -465 1471 -459 1 C3N
rlabel pdcontact 1457 -439 1461 -433 1 C3N
rlabel polycontact 1496 -434 1500 -430 1 C3N
rlabel ndcontact 1503 -440 1507 -436 1 C3
rlabel pdcontact 1503 -423 1507 -417 1 C3
rlabel ndcontact 1399 -451 1403 -447 1 gnd
rlabel pdcontact 1399 -433 1403 -427 1 vdd
rlabel nwell 1413 -425 1415 -423 1 vdd
rlabel polycontact 1400 -444 1404 -440 1 KP
rlabel ndcontact 1407 -450 1411 -446 1 KPK
rlabel pdcontact 1407 -433 1411 -427 1 KPK
rlabel polycontact 1468 -472 1472 -468 1 KPK
rlabel polycontact 1458 -394 1462 -390 1 KPK
rlabel pdcontact 1617 -300 1621 -288 1 vdd
rlabel pdcontact 1636 -282 1640 -270 1 vdd
rlabel pdcontact 1656 -268 1660 -256 1 vdd
rlabel polycontact 1641 -361 1645 -357 1 P2
rlabel polycontact 1637 -267 1641 -263 1 P2
rlabel pdcontact 1673 -248 1677 -236 1 vdd
rlabel polycontact 1674 -233 1678 -229 1 P3
rlabel polycontact 1657 -253 1661 -249 1 P1
rlabel polycontact 1641 -370 1645 -366 1 P1
rlabel polycontact 1641 -409 1645 -405 1 P3
rlabel polycontact 1618 -285 1622 -281 1 C1
rlabel polycontact 1641 -322 1645 -318 1 C1
rlabel pdcontact 1681 -245 1685 -239 1 AF
rlabel pdcontact 1664 -265 1668 -259 1 AF
rlabel pdcontact 1644 -278 1648 -272 1 AF
rlabel pdcontact 1625 -298 1629 -292 1 AF
rlabel ndcontact 1648 -333 1652 -327 1 AF
rlabel ndcontact 1640 -333 1644 -327 1 LO
rlabel ndcontact 1640 -354 1644 -348 1 LO
rlabel ndcontact 1648 -352 1652 -346 1 VE
rlabel ndcontact 1648 -380 1652 -374 1 VE
rlabel ndcontact 1640 -380 1644 -374 1 GA
rlabel ndcontact 1640 -401 1644 -395 1 GA
rlabel ndcontact 1648 -399 1652 -393 1 gnd
rlabel nwell 1631 -242 1633 -240 1 vdd
rlabel nwell 1705 -399 1707 -397 1 vdd
rlabel pdcontact 1691 -407 1695 -401 1 vdd
rlabel ndcontact 1691 -425 1695 -421 1 gnd
rlabel polycontact 1692 -418 1696 -414 1 AF
rlabel ndcontact 1699 -424 1703 -420 1 AFF
rlabel pdcontact 1699 -407 1703 -401 1 AFF
rlabel pdcontact 1985 -271 1989 -259 1 vdd
rlabel ndcontact 2003 -327 2007 -323 1 gnd
rlabel ndcontact 1977 -333 1981 -329 1 gnd
rlabel m123contact 1960 -326 1965 -321 1 HQ
rlabel polycontact 1978 -325 1982 -321 1 HQ
rlabel m123contact 1960 -288 1964 -284 1 HQ
rlabel polycontact 1986 -288 1990 -284 1 HQ
rlabel pdcontact 1993 -268 1997 -262 1 I2
rlabel pdcontact 1993 -299 1997 -293 1 I2
rlabel pdcontact 1985 -301 1989 -295 1 OJ
rlabel ndcontact 1985 -334 1989 -328 1 OJ
rlabel ndcontact 1995 -327 1999 -321 1 OJ
rlabel nwell 2000 -258 2002 -256 1 vdd
rlabel ndcontact 2030 -310 2034 -306 1 gnd
rlabel pdcontact 2030 -292 2034 -286 1 vdd
rlabel nwell 2044 -284 2046 -282 1 vdd
rlabel polycontact 2031 -303 2035 -299 1 OJ
rlabel ndcontact 2038 -309 2042 -305 1 OK
rlabel pdcontact 2038 -292 2042 -286 1 OK
rlabel m2contact 2065 -325 2068 -321 1 OK
rlabel pdcontact 1858 -292 1862 -280 1 vdd
rlabel pdcontact 1877 -274 1881 -262 1 vdd
rlabel pdcontact 1897 -260 1901 -248 1 vdd
rlabel ndcontact 1881 -374 1885 -365 1 gnd
rlabel polycontact 1898 -245 1902 -241 1 P3
rlabel polycontact 1882 -362 1886 -358 1 P3
rlabel polycontact 1882 -353 1886 -349 1 P2
rlabel polycontact 1878 -259 1882 -255 1 P2
rlabel polycontact 1859 -277 1863 -273 1 G1
rlabel polycontact 1882 -314 1886 -310 1 G1
rlabel ndcontact 1889 -371 1893 -367 1 AW
rlabel ndcontact 1889 -343 1893 -339 1 AW
rlabel ndcontact 1881 -345 1885 -341 1 NT
rlabel ndcontact 1881 -324 1885 -320 1 NT
rlabel ndcontact 1889 -324 1893 -320 1 LT
rlabel pdcontact 1866 -289 1870 -285 1 LT
rlabel pdcontact 1885 -269 1889 -265 1 LT
rlabel pdcontact 1905 -256 1909 -252 1 LT
rlabel nwell 1912 -245 1914 -243 1 vdd
rlabel ndcontact 1931 -313 1935 -309 1 gnd
rlabel pdcontact 1931 -295 1935 -289 1 vdd
rlabel nwell 1945 -287 1947 -285 1 vdd
rlabel polycontact 1932 -306 1936 -302 1 LT
rlabel ndcontact 1939 -312 1943 -308 1 6R
rlabel pdcontact 1939 -295 1943 -289 1 6R
rlabel polycontact 1996 -334 2000 -330 1 6R
rlabel polycontact 1986 -256 1990 -252 1 6R
rlabel pdcontact 2097 -271 2101 -259 1 vdd
rlabel ndcontact 2115 -327 2119 -323 1 gnd
rlabel ndcontact 2089 -333 2093 -329 1 gnd
rlabel pdcontact 2105 -268 2109 -262 1 I3
rlabel pdcontact 2105 -299 2109 -293 1 I3
rlabel nwell 2112 -256 2114 -254 1 vdd
rlabel ndcontact 2136 -307 2140 -303 1 gnd
rlabel pdcontact 2136 -289 2140 -283 1 vdd
rlabel nwell 2150 -281 2152 -279 1 vdd
rlabel ndcontact 2097 -334 2101 -328 1 C4N
rlabel ndcontact 2107 -327 2111 -321 1 C4N
rlabel pdcontact 2097 -301 2101 -295 1 C4N
rlabel polycontact 2137 -300 2141 -296 1 C4N
rlabel ndcontact 2144 -306 2148 -302 1 C4
rlabel pdcontact 2144 -289 2148 -283 1 C4
rlabel polycontact 2090 -325 2094 -321 1 OK
rlabel polycontact 2098 -256 2102 -252 1 OK
rlabel polycontact 2108 -334 2112 -330 1 AFF
rlabel polycontact 2098 -288 2102 -284 1 AFF
rlabel ndcontact 1737 -354 1741 -348 1 L34
rlabel pdcontact 1736 -303 1740 -297 1 L34
rlabel pdcontact 1775 -303 1779 -297 1 L34
rlabel ndcontact 1768 -341 1772 -335 1 L34
rlabel polycontact 1798 -332 1802 -328 1 L34
rlabel polycontact 1738 -361 1742 -357 1 G3
<< end >>
