.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd
.param width_P=2*width_N
.param width_N=3*LAMBDA

Vdd	vdd	gnd	'SUPPLY'
VX1 p1 gnd 1.8
VX2 c1 gnd pulse 0 1.8 0ns 100ps 100ps 10ns 20ns
VX4 p3 gnd 1.8
VX11 c3 gnd pulse 0 1.8 0ns 100ps 100ps 10ns 20ns
VX21 p2 gnd 1.8
VX31 c2 gnd pulse 0 1.8 0ns 100ps 100ps 10ns 20ns
VX41 p0 gnd 0
VX0 c0 gnd pulse 0 1.8 0ns 100ps 100ps 15ns 30ns

* SPICE3 file created from sum.ext - technology: scmos

.option scale=90n

M1000 S2 S2N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1001 C1N1 C1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1002 S0N C0N1 P0N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1003 C3N1 C3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1004 P1N1 P1 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1005 S2N C2N1 P2N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1006 S0 S0N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1007 P3N1 P3 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1008 P1N1 P1 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1009 S1N C1N1 P1N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1010 S0N C0 P0 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1011 S2N C2 P2 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1012 P3N1 P3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1013 S1N C1 P1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1014 C2N1 C2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1015 C1N1 C1 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1016 C3N1 C3 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1017 P2N1 P2 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1018 S0 S0N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1019 S1 S1N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1020 S3N C3N1 P3N1 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1021 P2N1 P2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1022 S3 S3N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1023 S1 S1N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1024 P0N1 P0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1025 S3N C3 P3 Gnd CMOSN w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1026 S3 S3N gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1027 C2N1 C2 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1028 P0N1 P0 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1029 S2 S2N vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1030 C0N1 C0 vdd vdd CMOSP w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1031 C0N1 C0 gnd Gnd CMOSN w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
C0 P1 C1 6.04e-19
C1 S2N m3_1218_n316# 1.12e-19
C2 vdd m2_723_n350# 0.00571f
C3 C0N1 gnd 0.072183f
C4 C3 C3N1 1.62e-19
C5 vdd C1N1 0.094864f
C6 P2 m3_1129_n299# 1.13e-19
C7 S0N m3_845_n320# 1.12e-19
C8 C0 m2_723_n350# 7.05e-19
C9 C2 gnd 0.056518f
C10 C3 vdd 0.043881f
C11 P0 m3_756_n303# 1.13e-19
C12 C0 gnd 0.056518f
C13 m2_1332_n348# m3_1332_n296# 4.06e-19
C14 P1N1 vdd 0.094864f
C15 P1 m3_946_n296# 1.13e-19
C16 S2 gnd 0.072183f
C17 C1 vdd 0.043881f
C18 P2 m2_1095_n346# 3.1e-19
C19 S3N gnd 0.080082f
C20 m2_1095_n346# m3_1129_n299# 0.007496f
C21 S0N gnd 0.080082f
C22 S0 vdd 0.094864f
C23 m2_723_n350# m3_756_n303# 0.007496f
C24 S3N C3 0.001447f
C25 S2N vdd 0.067556f
C26 P3 gnd 0.056518f
C27 vdd m3_1218_n316# 0.001729f
C28 P2 vdd 0.275061f
C29 S2N C2 0.001447f
C30 vdd m3_1129_n299# 0.001731f
C31 P2 C2 6.04e-19
C32 P3 C3 6.04e-19
C33 P1 vdd 0.275061f
C34 gnd m2_1300_n343# 0.002765f
C35 vdd m3_946_n296# 0.001731f
C36 P3N1 m2_1332_n348# 2.88e-19
C37 C0N1 m2_756_n355# 0.001081f
C38 P0 P0N1 1.62e-19
C39 S2N S2 1.62e-19
C40 S2 m3_1218_n316# 1.87e-19
C41 gnd m2_908_n343# 0.002765f
C42 vdd m2_756_n355# 0.004941f
C43 vdd m3_1421_n313# 0.001729f
C44 S0N S0 1.62e-19
C45 S1N S1 1.62e-19
C46 C2N1 gnd 0.072183f
C47 S1 m3_1035_n313# 1.87e-19
C48 vdd m2_1095_n346# 0.00571f
C49 C3 m2_1300_n343# 7.05e-19
C50 C0 m2_756_n355# 3.61e-19
C51 P3N1 gnd 0.072183f
C52 S1N m3_1035_n313# 1.12e-19
C53 vdd C3N1 0.094864f
C54 C2 m2_1095_n346# 7.05e-19
C55 P2N1 gnd 0.072183f
C56 vdd C0N1 0.094864f
C57 C1 m2_908_n343# 7.05e-19
C58 P0N1 gnd 0.072183f
C59 S3N m3_1421_n313# 1.12e-19
C60 C0 C0N1 1.62e-19
C61 S3 gnd 0.072183f
C62 C2 vdd 0.043881f
C63 m2_1129_n351# m3_1129_n299# 4.06e-19
C64 C0 vdd 0.043881f
C65 S1 gnd 0.072183f
C66 S3N C3N1 4.82e-19
C67 m2_756_n355# m3_756_n303# 4.06e-19
C68 P0 m2_723_n350# 3.1e-19
C69 S2N C2N1 4.82e-19
C70 S1N gnd 0.080082f
C71 S2 vdd 0.094864f
C72 S0N C0N1 4.82e-19
C73 S1N C1N1 4.82e-19
C74 P1 m2_908_n343# 3.1e-19
C75 S3N vdd 0.067556f
C76 P0 gnd 0.056518f
C77 m2_908_n343# m3_946_n296# 0.007496f
C78 S0N vdd 0.067556f
C79 vdd m3_1332_n296# 0.001731f
C80 P3 vdd 0.275061f
C81 P2 P2N1 1.62e-19
C82 vdd m3_756_n303# 0.001731f
C83 P2N1 m3_1129_n299# 3.33e-19
C84 S1N C1 0.001447f
C85 S0N C0 0.001447f
C86 vdd m2_1129_n351# 0.004941f
C87 C3 m2_1332_n348# 3.61e-19
C88 C1N1 m2_946_n348# 0.001081f
C89 gnd m2_723_n350# 0.002765f
C90 C2 m2_1129_n351# 3.61e-19
C91 vdd m2_1300_n343# 0.00571f
C92 P0N1 m2_756_n355# 2.88e-19
C93 C1N1 gnd 0.072183f
C94 P1N1 m2_946_n348# 2.88e-19
C95 S0 m3_845_n320# 1.87e-19
C96 vdd m2_908_n343# 0.00571f
C97 vdd C2N1 0.094864f
C98 C3 gnd 0.056518f
C99 C1 m2_946_n348# 3.61e-19
C100 S3 m3_1421_n313# 1.87e-19
C101 C2 C2N1 1.62e-19
C102 P3 m3_1332_n296# 1.13e-19
C103 P1N1 gnd 0.072183f
C104 vdd P3N1 0.094864f
C105 P2N1 vdd 0.094864f
C106 C1 gnd 0.056518f
C107 P0N1 vdd 0.094864f
C108 S0 gnd 0.072183f
C109 C1 C1N1 1.62e-19
C110 m2_1300_n343# m3_1332_n296# 0.007496f
C111 S2N gnd 0.080082f
C112 P3 m2_1300_n343# 3.1e-19
C113 S3 vdd 0.094864f
C114 m2_946_n348# m3_946_n296# 4.06e-19
C115 S1 vdd 0.094864f
C116 P2 gnd 0.056518f
C117 S1N vdd 0.067556f
C118 P1 gnd 0.056518f
C119 vdd m3_1035_n313# 0.001729f
C120 P3N1 m3_1332_n296# 3.33e-19
C121 C3N1 m2_1332_n348# 0.001081f
C122 P3 P3N1 1.62e-19
C123 P0 vdd 0.275061f
C124 vdd m3_845_n320# 0.001729f
C125 C2N1 m2_1129_n351# 0.001081f
C126 S3N S3 1.62e-19
C127 vdd m2_1332_n348# 0.004941f
C128 gnd m2_1095_n346# 0.002765f
C129 P1 P1N1 1.62e-19
C130 P0 C0 6.04e-19
C131 P2N1 m2_1129_n351# 2.88e-19
C132 gnd C3N1 0.072183f
C133 P0N1 m3_756_n303# 3.33e-19
C134 vdd m2_946_n348# 0.004941f
C135 P1N1 m3_946_n296# 3.33e-19
C136 m3_1421_n313# 0 0.016037f
C137 m3_1218_n316# 0 0.016037f
C138 m3_1035_n313# 0 0.016037f
C139 m3_1332_n296# 0 0.084889f
C140 m3_1129_n299# 0 0.084889f
C141 m3_845_n320# 0 0.016037f
C142 m3_756_n303# 0 0.084889f
C143 m3_946_n296# 0 0.084889f
C144 m2_1332_n348# 0 0.787321f
C145 m2_1129_n351# 0 0.787321f
C146 m2_756_n355# 0 0.787321f
C147 m2_946_n348# 0 0.787321f
C148 m2_1300_n343# 0 1.61989f
C149 m2_1095_n346# 0 1.642f
C150 m2_723_n350# 0 1.63095f
C151 m2_908_n343# 0 1.68623f
C152 C3N1 0 0.143763f 
C153 gnd 0 1.104016f 
C154 C2N1 0 0.143763f 
C155 C0N1 0 0.143763f 
C156 C1N1 0 0.143763f 
C157 P3N1 0 0.041372f 
C158 vdd 0 6.116681f 
C159 C3 0 0.281737f 
C160 P2N1 0 0.041372f 
C161 C2 0 0.281737f 
C162 P1N1 0 0.041372f 
C163 P0N1 0 0.041372f 
C164 C0 0 0.281737f 
C165 C1 0 0.281737f 
C166 S3 0 0.019328f 
C167 S2 0 0.019328f 
C168 S0 0 0.019328f 
C169 S1 0 0.019328f 
C170 S3N 0 0.320702f 
C171 S2N 0 0.320702f 
C172 S1N 0 0.320702f 
C173 S0N 0 0.320702f 
C174 P2 0 0.637785f 
C175 P0 0 0.634517f 
C176 P3 0 0.63125f 
C177 P1 0 0.650855f 



.tran 1n 80n 0n
.measure tran tpd_rise
+ TRIG v(b0) VAL='SUPPLY/2' RISE=1
+ TARG v(s3) VAL='SUPPLY/2' FALL=1
.measure tran tpd_fall
+ TRIG v(b0) VAL='SUPPLY/2' FALL=1
+ TARG v(s3) VAL='SUPPLY/2' RISE=1
.measure tran total_prop_delay param='(tpd_rise+tpd_fall)/2'
.control

run
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))
set curplottitle= harshita_2023102073

plot v(c0)+2 v(p0) v(s0)-2
plot v(p1)+2 v(c1) v(s1)-2
plot v(p2)+2 v(c2) v(s2)-2
plot v(p3)+2 v(c3) v(s3)-2

;plot v(c)

.endc