magic
tech scmos
timestamp 1731916657
<< nwell >>
rect 0 0 36 46
rect 70 14 104 49
rect 127 17 161 52
rect 183 23 208 53
<< ntransistor >>
rect 195 8 197 11
rect 142 -2 148 0
rect 85 -5 91 -3
rect 17 -14 20 -12
rect 142 -27 148 -25
rect 85 -30 91 -28
<< ptransistor >>
rect 141 38 147 40
rect 195 39 197 45
rect 84 35 90 37
rect 12 31 24 33
rect 12 13 24 15
<< ndiffusion >>
rect 194 8 195 11
rect 197 8 198 11
rect 89 -1 91 3
rect 146 2 148 6
rect 85 -3 91 -1
rect 142 0 148 2
rect 142 -3 148 -2
rect 85 -6 91 -5
rect 85 -10 86 -6
rect 90 -10 91 -6
rect 142 -7 143 -3
rect 147 -7 148 -3
rect 17 -12 20 -11
rect 17 -15 20 -14
rect 85 -26 86 -22
rect 90 -26 91 -22
rect 142 -23 143 -19
rect 147 -23 148 -19
rect 85 -28 91 -26
rect 142 -25 148 -23
rect 142 -28 148 -27
rect 85 -31 91 -30
rect 85 -35 86 -31
rect 90 -35 91 -31
rect 142 -32 143 -28
rect 147 -32 148 -28
<< pdiffusion >>
rect 84 38 85 42
rect 89 38 90 42
rect 141 41 142 45
rect 146 41 147 45
rect 12 34 16 38
rect 20 34 24 38
rect 84 37 90 38
rect 141 40 147 41
rect 194 39 195 45
rect 197 39 198 45
rect 141 37 147 38
rect 84 34 90 35
rect 12 33 24 34
rect 12 30 24 31
rect 84 30 85 34
rect 89 30 90 34
rect 141 33 142 37
rect 146 33 147 37
rect 12 26 16 30
rect 20 26 24 30
rect 12 16 16 20
rect 20 16 24 20
rect 12 15 24 16
rect 12 12 24 13
rect 12 8 16 12
rect 20 8 24 12
<< ndcontact >>
rect 190 7 194 11
rect 198 8 202 12
rect 85 -1 89 3
rect 142 2 146 6
rect 16 -11 20 -7
rect 86 -10 90 -6
rect 143 -7 147 -3
rect 16 -19 20 -15
rect 86 -26 90 -22
rect 143 -23 147 -19
rect 86 -35 90 -31
rect 143 -32 147 -28
<< pdcontact >>
rect 85 38 89 42
rect 142 41 146 45
rect 16 34 20 38
rect 190 39 194 45
rect 198 39 202 45
rect 85 30 89 34
rect 142 33 146 37
rect 16 26 20 30
rect 16 16 20 20
rect 16 8 20 12
<< polysilicon >>
rect 195 45 197 48
rect 135 38 141 40
rect 147 38 155 40
rect 78 35 84 37
rect 90 35 98 37
rect 5 31 12 33
rect 24 31 31 33
rect 5 13 12 15
rect 24 13 31 15
rect 195 11 197 39
rect 195 5 197 8
rect 134 -2 142 0
rect 148 -2 154 0
rect 77 -5 85 -3
rect 91 -5 97 -3
rect 5 -14 17 -12
rect 20 -14 31 -12
rect 134 -27 142 -25
rect 148 -27 154 -25
rect 77 -30 85 -28
rect 91 -30 97 -28
<< polycontact >>
rect 5 33 9 37
rect 74 34 78 38
rect 131 37 135 41
rect 5 15 9 19
rect 191 15 195 19
rect 73 -6 77 -2
rect 130 -3 134 1
rect 5 -12 9 -8
rect 73 -31 77 -27
rect 130 -28 134 -24
<< metal1 >>
rect 102 53 208 56
rect 33 52 208 53
rect 33 49 106 52
rect 127 51 208 52
rect 127 49 161 51
rect 33 48 37 49
rect 0 44 37 48
rect 70 47 106 49
rect 16 38 20 44
rect 85 42 89 47
rect 142 45 146 49
rect 190 45 194 51
rect 111 37 131 41
rect 16 20 20 26
rect 16 -2 20 8
rect 85 11 89 30
rect 111 11 115 37
rect 85 7 115 11
rect 85 3 89 7
rect 16 -6 73 -2
rect 16 -7 20 -6
rect 0 -23 34 -19
rect 30 -39 34 -23
rect 86 -22 90 -10
rect 111 -24 115 7
rect 142 14 146 33
rect 198 19 202 39
rect 177 15 191 19
rect 198 15 208 19
rect 177 14 181 15
rect 142 10 181 14
rect 198 12 202 15
rect 142 6 146 10
rect 190 -3 194 7
rect 143 -19 147 -7
rect 183 -7 208 -3
rect 111 -28 130 -24
rect 86 -39 90 -35
rect 143 -36 147 -32
rect 183 -36 187 -7
rect 129 -39 187 -36
rect 30 -40 187 -39
rect 30 -43 133 -40
<< labels >>
rlabel polycontact 5 -12 9 -8 1 D
rlabel polycontact 5 33 9 37 1 D
rlabel polycontact 5 15 9 19 1 clk
rlabel polycontact 73 -31 77 -27 1 clk
rlabel polycontact 74 34 78 38 1 clk
rlabel polycontact 130 -3 134 1 1 clk
rlabel metal1 204 15 208 19 7 Q
rlabel metal1 46 -6 52 -2 1 A
rlabel metal1 102 7 108 11 1 B
rlabel metal1 163 10 169 14 1 C
rlabel metal1 74 49 99 53 1 vdd
rlabel metal1 133 52 158 56 5 vdd
rlabel metal1 182 51 207 55 5 vdd
rlabel metal1 86 -19 90 -15 1 E
rlabel metal1 16 21 20 25 1 F
rlabel metal1 143 -16 147 -12 1 G
rlabel metal1 127 49 161 53 1 vdd
rlabel metal1 70 47 104 51 1 vdd
rlabel metal1 0 44 36 48 5 vdd
rlabel metal1 0 44 36 47 1 vdd
rlabel metal1 183 51 208 53 5 vdd
rlabel nwell 149 43 152 46 1 vdd
rlabel nwell 92 40 95 43 1 vdd
rlabel nwell 30 39 33 42 1 vdd
rlabel nwell 204 46 207 49 7 vdd
rlabel pdcontact 16 34 20 38 1 vdd
rlabel pdcontact 16 26 20 30 1 F
rlabel pdcontact 16 16 20 20 1 F
rlabel pdcontact 16 8 20 12 1 A
rlabel ndcontact 16 -11 20 -7 1 A
rlabel ndcontact 16 -19 20 -15 1 gnd
rlabel ndcontact 86 -35 90 -31 1 gnd
rlabel ndcontact 143 -32 147 -28 1 gnd
rlabel ndcontact 190 7 194 11 1 gnd
rlabel ndcontact 86 -26 90 -22 1 E
rlabel ndcontact 86 -10 90 -6 1 E
rlabel polycontact 73 -6 77 -2 1 A
rlabel ndcontact 85 -1 89 3 1 B
rlabel pdcontact 85 30 89 34 1 B
rlabel pdcontact 85 38 89 42 1 vdd
rlabel polycontact 130 -28 134 -24 1 B
rlabel ndcontact 143 -23 147 -19 1 G
rlabel ndcontact 143 -7 147 -3 1 G
rlabel ndcontact 142 2 146 6 1 C
rlabel pdcontact 142 33 146 37 1 C
rlabel pdcontact 142 41 146 45 1 vdd
rlabel polycontact 131 37 135 41 1 B
rlabel polycontact 191 15 195 19 1 C
rlabel pdcontact 190 39 194 45 1 vdd
rlabel pdcontact 198 39 202 45 1 Q
rlabel ndcontact 198 8 202 12 1 Q
<< end >>
