magic
tech scmos
timestamp 1732051476
<< nwell >>
rect 240 1271 276 1317
rect 310 1285 344 1320
rect 367 1288 401 1323
rect 423 1294 448 1324
rect 552 1250 576 1268
rect 641 1233 665 1251
rect 738 1247 762 1265
rect 827 1230 851 1248
rect 857 1220 893 1266
rect 927 1234 961 1269
rect 984 1237 1018 1272
rect 1040 1243 1065 1273
rect 1216 1239 1252 1285
rect 1258 1253 1292 1288
rect 1304 1256 1338 1291
rect 1344 1262 1369 1292
rect 1419 1270 1443 1288
rect 1508 1253 1532 1271
rect 1610 1267 1634 1285
rect 1699 1250 1723 1268
rect 1734 1240 1770 1286
rect 1776 1254 1810 1289
rect 1822 1257 1856 1292
rect 1862 1263 1887 1293
rect 1419 1218 1443 1236
rect 233 1162 269 1208
rect 303 1176 337 1211
rect 360 1179 394 1214
rect 416 1185 441 1215
rect 552 1198 576 1216
rect 1610 1215 1634 1233
rect 738 1195 762 1213
rect 657 1147 717 1181
rect 1239 1131 1275 1177
rect 1281 1145 1315 1180
rect 1327 1148 1361 1183
rect 1367 1154 1392 1184
rect 1414 1125 1474 1159
rect 389 1044 425 1090
rect 459 1058 493 1093
rect 516 1061 550 1096
rect 572 1067 597 1097
rect 798 1090 858 1124
rect 1469 1093 1493 1111
rect 1558 1093 1619 1155
rect 1715 1106 1784 1166
rect 1799 1106 1823 1124
rect 1625 1080 1649 1098
rect 1861 1097 1886 1154
rect 1895 1109 1919 1127
rect 658 1011 718 1045
rect 739 860 775 906
rect 786 874 820 909
rect 843 877 877 912
rect 899 883 924 913
rect 953 880 977 898
rect 1042 863 1066 881
rect 1114 877 1138 895
rect 1203 860 1227 878
rect 953 828 977 846
rect 1114 825 1138 843
rect 1248 836 1284 882
rect 1294 850 1328 885
rect 1351 853 1385 888
rect 1397 859 1422 889
rect 1661 790 1697 836
rect 1703 804 1737 839
rect 1749 807 1783 842
rect 1789 813 1814 843
rect 1841 810 1865 828
rect 1930 793 1954 811
rect 2101 807 2125 825
rect 2190 790 2214 808
rect 769 729 805 775
rect 811 743 845 778
rect 860 746 894 781
rect 903 752 928 782
rect 948 737 1008 771
rect 1003 705 1027 723
rect 1092 717 1153 779
rect 1841 758 1865 776
rect 2101 755 2125 773
rect 2225 770 2261 816
rect 2267 784 2301 819
rect 2313 787 2347 822
rect 2353 793 2378 823
rect 1159 704 1183 722
rect 1661 648 1697 694
rect 1703 662 1737 697
rect 1749 665 1783 700
rect 1789 671 1814 701
rect 1836 606 1896 640
rect 2019 620 2105 702
rect 2167 615 2228 677
rect 2295 628 2364 688
rect 2375 628 2399 646
rect 2234 602 2258 620
rect 2433 619 2458 676
rect 2479 619 2503 637
rect 2562 619 2587 676
rect 2597 619 2621 637
rect 2640 626 2676 672
rect 2682 640 2716 675
rect 2728 643 2762 678
rect 2768 649 2793 679
rect 1895 574 1919 592
rect 2107 516 2131 534
<< ntransistor >>
rect 435 1279 437 1282
rect 382 1269 388 1271
rect 325 1266 331 1268
rect 257 1257 260 1259
rect 382 1244 388 1246
rect 325 1241 331 1243
rect 622 1250 624 1256
rect 563 1239 565 1242
rect 808 1247 810 1253
rect 749 1236 751 1239
rect 652 1222 654 1225
rect 1489 1270 1491 1276
rect 1430 1259 1432 1262
rect 1680 1267 1682 1273
rect 1356 1247 1358 1250
rect 1621 1256 1623 1259
rect 1519 1242 1521 1245
rect 1874 1248 1876 1251
rect 1319 1237 1325 1239
rect 1710 1239 1712 1242
rect 1273 1234 1279 1236
rect 1052 1228 1054 1231
rect 838 1219 840 1222
rect 1233 1225 1236 1227
rect 1489 1229 1491 1235
rect 1837 1238 1843 1240
rect 1791 1235 1797 1237
rect 622 1209 624 1215
rect 999 1218 1005 1220
rect 942 1215 948 1217
rect 808 1206 810 1212
rect 1680 1226 1682 1232
rect 1751 1226 1754 1228
rect 1319 1212 1325 1214
rect 1273 1209 1279 1211
rect 874 1206 877 1208
rect 1430 1207 1432 1210
rect 1837 1213 1843 1215
rect 1791 1210 1797 1212
rect 1621 1204 1623 1207
rect 563 1187 565 1190
rect 999 1193 1005 1195
rect 942 1190 948 1192
rect 749 1184 751 1187
rect 428 1170 430 1173
rect 375 1160 381 1162
rect 318 1157 324 1159
rect 250 1148 253 1150
rect 1379 1139 1381 1142
rect 375 1135 381 1137
rect 318 1132 324 1134
rect 686 1120 688 1126
rect 1342 1129 1348 1131
rect 1296 1126 1302 1128
rect 1256 1117 1259 1119
rect 686 1094 688 1100
rect 1342 1104 1348 1106
rect 1296 1101 1302 1103
rect 1443 1098 1445 1104
rect 1810 1095 1812 1098
rect 1906 1098 1908 1101
rect 1480 1082 1482 1085
rect 1443 1072 1445 1078
rect 1754 1081 1756 1090
rect 1883 1080 1885 1086
rect 1865 1073 1867 1079
rect 827 1063 829 1069
rect 1599 1066 1601 1072
rect 1636 1069 1638 1072
rect 1754 1061 1756 1070
rect 584 1052 586 1055
rect 1576 1053 1578 1059
rect 531 1042 537 1044
rect 474 1039 480 1041
rect 827 1037 829 1043
rect 1599 1040 1601 1046
rect 406 1030 409 1032
rect 1754 1033 1756 1042
rect 531 1017 537 1019
rect 474 1014 480 1016
rect 687 984 689 990
rect 687 958 689 964
rect 1023 880 1025 886
rect 911 868 913 871
rect 964 869 966 872
rect 1184 877 1186 883
rect 858 858 864 860
rect 801 855 807 857
rect 1125 866 1127 869
rect 1053 852 1055 855
rect 1214 849 1216 852
rect 756 846 759 848
rect 858 833 864 835
rect 1023 839 1025 845
rect 1409 844 1411 847
rect 801 830 807 832
rect 1184 836 1186 842
rect 1366 834 1372 836
rect 1309 831 1315 833
rect 964 817 966 820
rect 1265 822 1268 824
rect 1125 814 1127 817
rect 1366 809 1372 811
rect 1309 806 1315 808
rect 1911 810 1913 816
rect 1801 798 1803 801
rect 1852 799 1854 802
rect 2171 807 2173 813
rect 1764 788 1770 790
rect 1718 785 1724 787
rect 2112 796 2114 799
rect 1941 782 1943 785
rect 2201 779 2203 782
rect 1678 776 1681 778
rect 2365 778 2367 781
rect 1764 763 1770 765
rect 1911 769 1913 775
rect 1718 760 1724 762
rect 2171 766 2173 772
rect 2328 768 2334 770
rect 2282 765 2288 767
rect 2242 756 2245 758
rect 1852 747 1854 750
rect 915 737 917 740
rect 2112 744 2114 747
rect 2328 743 2334 745
rect 2282 740 2288 742
rect 875 727 881 729
rect 826 724 832 726
rect 786 715 789 717
rect 977 710 979 716
rect 875 702 881 704
rect 826 699 832 701
rect 1014 694 1016 697
rect 1133 690 1135 696
rect 1170 693 1172 696
rect 977 684 979 690
rect 1110 677 1112 683
rect 1133 664 1135 670
rect 1801 656 1803 659
rect 1764 646 1770 648
rect 1718 643 1724 645
rect 1678 634 1681 636
rect 1764 621 1770 623
rect 1718 618 1724 620
rect 2780 634 2782 637
rect 2386 617 2388 620
rect 2058 595 2060 604
rect 2334 603 2336 612
rect 2455 602 2457 608
rect 2490 608 2492 611
rect 2743 624 2749 626
rect 2697 621 2703 623
rect 2657 612 2660 614
rect 2437 595 2439 601
rect 2584 602 2586 608
rect 2608 608 2610 611
rect 2566 595 2568 601
rect 2743 599 2749 601
rect 2697 596 2703 598
rect 2208 588 2210 594
rect 2245 591 2247 594
rect 1865 579 1867 585
rect 2058 575 2060 584
rect 2334 583 2336 592
rect 2185 575 2187 581
rect 1906 563 1908 566
rect 1865 553 1867 559
rect 2208 562 2210 568
rect 2058 547 2060 556
rect 2334 555 2336 564
rect 2058 527 2060 536
rect 2118 505 2120 508
<< ptransistor >>
rect 381 1309 387 1311
rect 435 1310 437 1316
rect 324 1306 330 1308
rect 252 1302 264 1304
rect 252 1284 264 1286
rect 1318 1277 1324 1279
rect 1356 1278 1358 1284
rect 1272 1274 1278 1276
rect 1228 1270 1240 1272
rect 563 1256 565 1262
rect 749 1253 751 1259
rect 998 1258 1004 1260
rect 1052 1259 1054 1265
rect 941 1255 947 1257
rect 652 1239 654 1245
rect 869 1251 881 1253
rect 838 1236 840 1242
rect 869 1233 881 1235
rect 1228 1252 1240 1254
rect 1430 1276 1432 1282
rect 1621 1273 1623 1279
rect 1836 1278 1842 1280
rect 1874 1279 1876 1285
rect 1790 1275 1796 1277
rect 1519 1259 1521 1265
rect 1746 1271 1758 1273
rect 1710 1256 1712 1262
rect 1746 1253 1758 1255
rect 1430 1224 1432 1230
rect 374 1200 380 1202
rect 428 1201 430 1207
rect 563 1204 565 1210
rect 317 1197 323 1199
rect 245 1193 257 1195
rect 245 1175 257 1177
rect 749 1201 751 1207
rect 1621 1221 1623 1227
rect 678 1169 680 1175
rect 1341 1169 1347 1171
rect 1379 1170 1381 1176
rect 1295 1166 1301 1168
rect 1251 1162 1263 1164
rect 704 1153 706 1159
rect 1251 1144 1263 1146
rect 1435 1147 1437 1153
rect 1461 1131 1463 1137
rect 1583 1135 1585 1147
rect 1770 1147 1772 1159
rect 1750 1133 1752 1145
rect 1873 1136 1875 1148
rect 819 1112 821 1118
rect 1731 1115 1733 1127
rect 845 1096 847 1102
rect 1480 1099 1482 1105
rect 1575 1101 1577 1113
rect 1606 1101 1608 1113
rect 1810 1112 1812 1118
rect 530 1082 536 1084
rect 584 1083 586 1089
rect 1873 1104 1875 1116
rect 1906 1115 1908 1121
rect 1636 1086 1638 1092
rect 473 1079 479 1081
rect 401 1075 413 1077
rect 401 1057 413 1059
rect 679 1033 681 1039
rect 705 1017 707 1023
rect 857 898 863 900
rect 911 899 913 905
rect 800 895 806 897
rect 751 891 763 893
rect 751 873 763 875
rect 964 886 966 892
rect 1125 883 1127 889
rect 1053 869 1055 875
rect 1214 866 1216 872
rect 1365 874 1371 876
rect 1409 875 1411 881
rect 1308 871 1314 873
rect 1260 867 1272 869
rect 1260 849 1272 851
rect 964 834 966 840
rect 1125 831 1127 837
rect 1763 828 1769 830
rect 1801 829 1803 835
rect 1717 825 1723 827
rect 1673 821 1685 823
rect 1673 803 1685 805
rect 1852 816 1854 822
rect 2112 813 2114 819
rect 1941 799 1943 805
rect 2327 808 2333 810
rect 2365 809 2367 815
rect 2281 805 2287 807
rect 2201 796 2203 802
rect 2237 801 2249 803
rect 2237 783 2249 785
rect 874 767 880 769
rect 915 768 917 774
rect 825 764 831 766
rect 781 760 793 762
rect 781 742 793 744
rect 969 759 971 765
rect 1117 759 1119 771
rect 1852 764 1854 770
rect 2112 761 2114 767
rect 995 743 997 749
rect 1109 725 1111 737
rect 1140 725 1142 737
rect 1014 711 1016 717
rect 1170 710 1172 716
rect 1763 686 1769 688
rect 1801 687 1803 693
rect 1717 683 1723 685
rect 1673 679 1685 681
rect 1673 661 1685 663
rect 2091 681 2093 693
rect 2074 661 2076 673
rect 2054 647 2056 659
rect 2192 657 2194 669
rect 2350 669 2352 681
rect 2330 655 2332 667
rect 2445 658 2447 670
rect 2574 658 2576 670
rect 2742 664 2748 666
rect 2780 665 2782 671
rect 2696 661 2702 663
rect 2652 657 2664 659
rect 1857 628 1859 634
rect 2035 629 2037 641
rect 2311 637 2313 649
rect 2184 623 2186 635
rect 2215 623 2217 635
rect 2386 634 2388 640
rect 2652 639 2664 641
rect 1883 612 1885 618
rect 2445 626 2447 638
rect 2490 625 2492 631
rect 2574 626 2576 638
rect 2245 608 2247 614
rect 2608 625 2610 631
rect 1906 580 1908 586
rect 2118 522 2120 528
<< ndiffusion >>
rect 434 1279 435 1282
rect 437 1279 438 1282
rect 329 1270 331 1274
rect 386 1273 388 1277
rect 325 1268 331 1270
rect 382 1271 388 1273
rect 382 1268 388 1269
rect 325 1265 331 1266
rect 325 1261 326 1265
rect 330 1261 331 1265
rect 382 1264 383 1268
rect 387 1264 388 1268
rect 257 1259 260 1260
rect 257 1256 260 1257
rect 325 1245 326 1249
rect 330 1245 331 1249
rect 382 1248 383 1252
rect 387 1248 388 1252
rect 325 1243 331 1245
rect 382 1246 388 1248
rect 382 1243 388 1244
rect 325 1240 331 1241
rect 325 1236 326 1240
rect 330 1236 331 1240
rect 382 1239 383 1243
rect 387 1239 388 1243
rect 617 1250 622 1256
rect 624 1250 630 1256
rect 562 1239 563 1242
rect 565 1239 566 1242
rect 803 1247 808 1253
rect 810 1247 816 1253
rect 748 1236 749 1239
rect 751 1236 752 1239
rect 651 1222 652 1225
rect 654 1222 655 1225
rect 1484 1270 1489 1276
rect 1491 1270 1497 1276
rect 1429 1259 1430 1262
rect 1432 1259 1433 1262
rect 1675 1267 1680 1273
rect 1682 1267 1688 1273
rect 1355 1247 1356 1250
rect 1358 1247 1359 1250
rect 1277 1238 1279 1242
rect 1323 1241 1325 1245
rect 1620 1256 1621 1259
rect 1623 1256 1624 1259
rect 1518 1242 1519 1245
rect 1521 1242 1522 1245
rect 1873 1248 1874 1251
rect 1876 1248 1877 1251
rect 1273 1236 1279 1238
rect 1319 1239 1325 1241
rect 1709 1239 1710 1242
rect 1712 1239 1713 1242
rect 1795 1239 1797 1243
rect 1841 1242 1843 1246
rect 1319 1236 1325 1237
rect 1273 1233 1279 1234
rect 1051 1228 1052 1231
rect 1054 1228 1055 1231
rect 837 1219 838 1222
rect 840 1219 841 1222
rect 946 1219 948 1223
rect 1003 1222 1005 1226
rect 1273 1229 1274 1233
rect 1278 1229 1279 1233
rect 1319 1232 1320 1236
rect 1324 1232 1325 1236
rect 1233 1227 1236 1228
rect 1233 1224 1236 1225
rect 1485 1229 1489 1235
rect 1491 1229 1497 1235
rect 1791 1237 1797 1239
rect 1837 1240 1843 1242
rect 1837 1237 1843 1238
rect 1791 1234 1797 1235
rect 618 1209 622 1215
rect 624 1209 630 1215
rect 942 1217 948 1219
rect 999 1220 1005 1222
rect 999 1217 1005 1218
rect 942 1214 948 1215
rect 804 1206 808 1212
rect 810 1206 816 1212
rect 942 1210 943 1214
rect 947 1210 948 1214
rect 999 1213 1000 1217
rect 1004 1213 1005 1217
rect 1273 1213 1274 1217
rect 1278 1213 1279 1217
rect 1319 1216 1320 1220
rect 1324 1216 1325 1220
rect 1676 1226 1680 1232
rect 1682 1226 1688 1232
rect 1791 1230 1792 1234
rect 1796 1230 1797 1234
rect 1837 1233 1838 1237
rect 1842 1233 1843 1237
rect 1751 1228 1754 1229
rect 874 1208 877 1209
rect 1273 1211 1279 1213
rect 1319 1214 1325 1216
rect 1751 1225 1754 1226
rect 1319 1211 1325 1212
rect 1273 1208 1279 1209
rect 874 1205 877 1206
rect 1273 1204 1274 1208
rect 1278 1204 1279 1208
rect 1319 1207 1320 1211
rect 1324 1207 1325 1211
rect 1429 1207 1430 1210
rect 1432 1207 1433 1210
rect 1791 1214 1792 1218
rect 1796 1214 1797 1218
rect 1837 1217 1838 1221
rect 1842 1217 1843 1221
rect 1791 1212 1797 1214
rect 1837 1215 1843 1217
rect 1837 1212 1843 1213
rect 1791 1209 1797 1210
rect 1620 1204 1621 1207
rect 1623 1204 1624 1207
rect 1791 1205 1792 1209
rect 1796 1205 1797 1209
rect 1837 1208 1838 1212
rect 1842 1208 1843 1212
rect 562 1187 563 1190
rect 565 1187 566 1190
rect 942 1194 943 1198
rect 947 1194 948 1198
rect 999 1197 1000 1201
rect 1004 1197 1005 1201
rect 942 1192 948 1194
rect 999 1195 1005 1197
rect 999 1192 1005 1193
rect 942 1189 948 1190
rect 748 1184 749 1187
rect 751 1184 752 1187
rect 942 1185 943 1189
rect 947 1185 948 1189
rect 999 1188 1000 1192
rect 1004 1188 1005 1192
rect 427 1170 428 1173
rect 430 1170 431 1173
rect 322 1161 324 1165
rect 379 1164 381 1168
rect 318 1159 324 1161
rect 375 1162 381 1164
rect 375 1159 381 1160
rect 318 1156 324 1157
rect 318 1152 319 1156
rect 323 1152 324 1156
rect 375 1155 376 1159
rect 380 1155 381 1159
rect 250 1150 253 1151
rect 250 1147 253 1148
rect 318 1136 319 1140
rect 323 1136 324 1140
rect 375 1139 376 1143
rect 380 1139 381 1143
rect 318 1134 324 1136
rect 375 1137 381 1139
rect 1378 1139 1379 1142
rect 1381 1139 1382 1142
rect 375 1134 381 1135
rect 318 1131 324 1132
rect 318 1127 319 1131
rect 323 1127 324 1131
rect 375 1130 376 1134
rect 380 1130 381 1134
rect 1300 1130 1302 1134
rect 1346 1133 1348 1137
rect 685 1120 686 1126
rect 688 1120 689 1126
rect 1296 1128 1302 1130
rect 1342 1131 1348 1133
rect 1342 1128 1348 1129
rect 1296 1125 1302 1126
rect 1296 1121 1297 1125
rect 1301 1121 1302 1125
rect 1342 1124 1343 1128
rect 1347 1124 1348 1128
rect 1256 1119 1259 1120
rect 1256 1116 1259 1117
rect 1296 1105 1297 1109
rect 1301 1105 1302 1109
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 685 1094 686 1100
rect 688 1094 689 1100
rect 1296 1103 1302 1105
rect 1342 1106 1348 1108
rect 1342 1103 1348 1104
rect 1296 1100 1302 1101
rect 1296 1096 1297 1100
rect 1301 1096 1302 1100
rect 1342 1099 1343 1103
rect 1347 1099 1348 1103
rect 1442 1098 1443 1104
rect 1445 1098 1446 1104
rect 1809 1095 1810 1098
rect 1812 1095 1813 1098
rect 1905 1098 1906 1101
rect 1908 1098 1909 1101
rect 1479 1082 1480 1085
rect 1482 1082 1483 1085
rect 1442 1072 1443 1078
rect 1445 1072 1446 1078
rect 1753 1081 1754 1090
rect 1756 1081 1757 1090
rect 1882 1080 1883 1086
rect 1885 1080 1886 1086
rect 1864 1073 1865 1079
rect 1867 1073 1868 1079
rect 826 1063 827 1069
rect 829 1063 830 1069
rect 1598 1066 1599 1072
rect 1601 1066 1602 1072
rect 1635 1069 1636 1072
rect 1638 1069 1639 1072
rect 1753 1061 1754 1070
rect 1756 1061 1757 1070
rect 583 1052 584 1055
rect 586 1052 587 1055
rect 1575 1053 1576 1059
rect 1578 1053 1579 1059
rect 478 1043 480 1047
rect 535 1046 537 1050
rect 474 1041 480 1043
rect 531 1044 537 1046
rect 531 1041 537 1042
rect 474 1038 480 1039
rect 474 1034 475 1038
rect 479 1034 480 1038
rect 531 1037 532 1041
rect 536 1037 537 1041
rect 826 1037 827 1043
rect 829 1037 830 1043
rect 1598 1040 1599 1046
rect 1601 1040 1602 1046
rect 406 1032 409 1033
rect 406 1029 409 1030
rect 1753 1033 1754 1042
rect 1756 1033 1757 1042
rect 474 1018 475 1022
rect 479 1018 480 1022
rect 531 1021 532 1025
rect 536 1021 537 1025
rect 474 1016 480 1018
rect 531 1019 537 1021
rect 531 1016 537 1017
rect 474 1013 480 1014
rect 474 1009 475 1013
rect 479 1009 480 1013
rect 531 1012 532 1016
rect 536 1012 537 1016
rect 686 984 687 990
rect 689 984 690 990
rect 686 958 687 964
rect 689 958 690 964
rect 1018 880 1023 886
rect 1025 880 1031 886
rect 910 868 911 871
rect 913 868 914 871
rect 963 869 964 872
rect 966 869 967 872
rect 1179 877 1184 883
rect 1186 877 1192 883
rect 805 859 807 863
rect 862 862 864 866
rect 801 857 807 859
rect 858 860 864 862
rect 858 857 864 858
rect 801 854 807 855
rect 801 850 802 854
rect 806 850 807 854
rect 858 853 859 857
rect 863 853 864 857
rect 1124 866 1125 869
rect 1127 866 1128 869
rect 1052 852 1053 855
rect 1055 852 1056 855
rect 756 848 759 849
rect 1213 849 1214 852
rect 1216 849 1217 852
rect 756 845 759 846
rect 801 834 802 838
rect 806 834 807 838
rect 858 837 859 841
rect 863 837 864 841
rect 801 832 807 834
rect 858 835 864 837
rect 1019 839 1023 845
rect 1025 839 1031 845
rect 1408 844 1409 847
rect 1411 844 1412 847
rect 858 832 864 833
rect 801 829 807 830
rect 801 825 802 829
rect 806 825 807 829
rect 858 828 859 832
rect 863 828 864 832
rect 1180 836 1184 842
rect 1186 836 1192 842
rect 1313 835 1315 839
rect 1370 838 1372 842
rect 1309 833 1315 835
rect 1366 836 1372 838
rect 1366 833 1372 834
rect 1309 830 1315 831
rect 963 817 964 820
rect 966 817 967 820
rect 1309 826 1310 830
rect 1314 826 1315 830
rect 1366 829 1367 833
rect 1371 829 1372 833
rect 1265 824 1268 825
rect 1265 821 1268 822
rect 1124 814 1125 817
rect 1127 814 1128 817
rect 1309 810 1310 814
rect 1314 810 1315 814
rect 1366 813 1367 817
rect 1371 813 1372 817
rect 1309 808 1315 810
rect 1366 811 1372 813
rect 1366 808 1372 809
rect 1309 805 1315 806
rect 1309 801 1310 805
rect 1314 801 1315 805
rect 1366 804 1367 808
rect 1371 804 1372 808
rect 1906 810 1911 816
rect 1913 810 1919 816
rect 1800 798 1801 801
rect 1803 798 1804 801
rect 1851 799 1852 802
rect 1854 799 1855 802
rect 2166 807 2171 813
rect 2173 807 2179 813
rect 1722 789 1724 793
rect 1768 792 1770 796
rect 1718 787 1724 789
rect 1764 790 1770 792
rect 1764 787 1770 788
rect 1718 784 1724 785
rect 1718 780 1719 784
rect 1723 780 1724 784
rect 1764 783 1765 787
rect 1769 783 1770 787
rect 2111 796 2112 799
rect 2114 796 2115 799
rect 1940 782 1941 785
rect 1943 782 1944 785
rect 1678 778 1681 779
rect 2200 779 2201 782
rect 2203 779 2204 782
rect 1678 775 1681 776
rect 2364 778 2365 781
rect 2367 778 2368 781
rect 1718 764 1719 768
rect 1723 764 1724 768
rect 1764 767 1765 771
rect 1769 767 1770 771
rect 1718 762 1724 764
rect 1764 765 1770 767
rect 1907 769 1911 775
rect 1913 769 1919 775
rect 1764 762 1770 763
rect 1718 759 1724 760
rect 1718 755 1719 759
rect 1723 755 1724 759
rect 1764 758 1765 762
rect 1769 758 1770 762
rect 2167 766 2171 772
rect 2173 766 2179 772
rect 2286 769 2288 773
rect 2332 772 2334 776
rect 2282 767 2288 769
rect 2328 770 2334 772
rect 2328 767 2334 768
rect 2282 764 2288 765
rect 2282 760 2283 764
rect 2287 760 2288 764
rect 2328 763 2329 767
rect 2333 763 2334 767
rect 2242 758 2245 759
rect 2242 755 2245 756
rect 1851 747 1852 750
rect 1854 747 1855 750
rect 914 737 915 740
rect 917 737 918 740
rect 2111 744 2112 747
rect 2114 744 2115 747
rect 2282 744 2283 748
rect 2287 744 2288 748
rect 2328 747 2329 751
rect 2333 747 2334 751
rect 2282 742 2288 744
rect 2328 745 2334 747
rect 2328 742 2334 743
rect 2282 739 2288 740
rect 830 728 832 732
rect 879 731 881 735
rect 826 726 832 728
rect 875 729 881 731
rect 875 726 881 727
rect 826 723 832 724
rect 826 719 827 723
rect 831 719 832 723
rect 875 722 876 726
rect 880 722 881 726
rect 2282 735 2283 739
rect 2287 735 2288 739
rect 2328 738 2329 742
rect 2333 738 2334 742
rect 786 717 789 718
rect 786 714 789 715
rect 976 710 977 716
rect 979 710 980 716
rect 826 703 827 707
rect 831 703 832 707
rect 875 706 876 710
rect 880 706 881 710
rect 826 701 832 703
rect 875 704 881 706
rect 875 701 881 702
rect 826 698 832 699
rect 826 694 827 698
rect 831 694 832 698
rect 875 697 876 701
rect 880 697 881 701
rect 1013 694 1014 697
rect 1016 694 1017 697
rect 1132 690 1133 696
rect 1135 690 1136 696
rect 1169 693 1170 696
rect 1172 693 1173 696
rect 976 684 977 690
rect 979 684 980 690
rect 1109 677 1110 683
rect 1112 677 1113 683
rect 1132 664 1133 670
rect 1135 664 1136 670
rect 1800 656 1801 659
rect 1803 656 1804 659
rect 1722 647 1724 651
rect 1768 650 1770 654
rect 1718 645 1724 647
rect 1764 648 1770 650
rect 1764 645 1770 646
rect 1718 642 1724 643
rect 1718 638 1719 642
rect 1723 638 1724 642
rect 1764 641 1765 645
rect 1769 641 1770 645
rect 1678 636 1681 637
rect 1678 633 1681 634
rect 1718 622 1719 626
rect 1723 622 1724 626
rect 1764 625 1765 629
rect 1769 625 1770 629
rect 1718 620 1724 622
rect 1764 623 1770 625
rect 1764 620 1770 621
rect 1718 617 1724 618
rect 1718 613 1719 617
rect 1723 613 1724 617
rect 1764 616 1765 620
rect 1769 616 1770 620
rect 2779 634 2780 637
rect 2782 634 2783 637
rect 2385 617 2386 620
rect 2388 617 2389 620
rect 2057 595 2058 604
rect 2060 595 2061 604
rect 2333 603 2334 612
rect 2336 603 2337 612
rect 2701 625 2703 629
rect 2747 628 2749 632
rect 2454 602 2455 608
rect 2457 602 2458 608
rect 2489 608 2490 611
rect 2492 608 2493 611
rect 2697 623 2703 625
rect 2743 626 2749 628
rect 2743 623 2749 624
rect 2697 620 2703 621
rect 2697 616 2698 620
rect 2702 616 2703 620
rect 2743 619 2744 623
rect 2748 619 2749 623
rect 2657 614 2660 615
rect 2436 595 2437 601
rect 2439 595 2440 601
rect 2583 602 2584 608
rect 2586 602 2587 608
rect 2607 608 2608 611
rect 2610 608 2611 611
rect 2657 611 2660 612
rect 2565 595 2566 601
rect 2568 595 2569 601
rect 2697 600 2698 604
rect 2702 600 2703 604
rect 2743 603 2744 607
rect 2748 603 2749 607
rect 2697 598 2703 600
rect 2743 601 2749 603
rect 2743 598 2749 599
rect 2697 595 2703 596
rect 2207 588 2208 594
rect 2210 588 2211 594
rect 2244 591 2245 594
rect 2247 591 2248 594
rect 1864 579 1865 585
rect 1867 579 1868 585
rect 2057 575 2058 584
rect 2060 575 2061 584
rect 2333 583 2334 592
rect 2336 583 2337 592
rect 2697 591 2698 595
rect 2702 591 2703 595
rect 2743 594 2744 598
rect 2748 594 2749 598
rect 2184 575 2185 581
rect 2187 575 2188 581
rect 1905 563 1906 566
rect 1908 563 1909 566
rect 1864 553 1865 559
rect 1867 553 1868 559
rect 2207 562 2208 568
rect 2210 562 2211 568
rect 2057 547 2058 556
rect 2060 547 2061 556
rect 2333 555 2334 564
rect 2336 555 2337 564
rect 2057 527 2058 536
rect 2060 527 2061 536
rect 2117 505 2118 508
rect 2120 505 2121 508
<< pdiffusion >>
rect 324 1309 325 1313
rect 329 1309 330 1313
rect 381 1312 382 1316
rect 386 1312 387 1316
rect 252 1305 256 1309
rect 260 1305 264 1309
rect 324 1308 330 1309
rect 381 1311 387 1312
rect 434 1310 435 1316
rect 437 1310 438 1316
rect 381 1308 387 1309
rect 324 1305 330 1306
rect 252 1304 264 1305
rect 252 1301 264 1302
rect 324 1301 325 1305
rect 329 1301 330 1305
rect 381 1304 382 1308
rect 386 1304 387 1308
rect 252 1297 256 1301
rect 260 1297 264 1301
rect 252 1287 256 1291
rect 260 1287 264 1291
rect 252 1286 264 1287
rect 252 1283 264 1284
rect 252 1279 256 1283
rect 260 1279 264 1283
rect 1272 1277 1273 1281
rect 1277 1277 1278 1281
rect 1318 1280 1319 1284
rect 1323 1280 1324 1284
rect 1228 1273 1232 1277
rect 1236 1273 1240 1277
rect 1272 1276 1278 1277
rect 1318 1279 1324 1280
rect 1355 1278 1356 1284
rect 1358 1278 1359 1284
rect 1318 1276 1324 1277
rect 1272 1273 1278 1274
rect 1228 1272 1240 1273
rect 1228 1269 1240 1270
rect 1272 1269 1273 1273
rect 1277 1269 1278 1273
rect 1318 1272 1319 1276
rect 1323 1272 1324 1276
rect 1228 1265 1232 1269
rect 1236 1265 1240 1269
rect 562 1256 563 1262
rect 565 1256 566 1262
rect 748 1253 749 1259
rect 751 1253 752 1259
rect 941 1258 942 1262
rect 946 1258 947 1262
rect 998 1261 999 1265
rect 1003 1261 1004 1265
rect 869 1254 873 1258
rect 877 1254 881 1258
rect 941 1257 947 1258
rect 998 1260 1004 1261
rect 1051 1259 1052 1265
rect 1054 1259 1055 1265
rect 998 1257 1004 1258
rect 941 1254 947 1255
rect 869 1253 881 1254
rect 651 1239 652 1245
rect 654 1239 655 1245
rect 869 1250 881 1251
rect 941 1250 942 1254
rect 946 1250 947 1254
rect 998 1253 999 1257
rect 1003 1253 1004 1257
rect 869 1246 873 1250
rect 877 1246 881 1250
rect 837 1236 838 1242
rect 840 1236 841 1242
rect 869 1236 873 1240
rect 877 1236 881 1240
rect 869 1235 881 1236
rect 869 1232 881 1233
rect 869 1228 873 1232
rect 877 1228 881 1232
rect 1228 1255 1232 1259
rect 1236 1255 1240 1259
rect 1228 1254 1240 1255
rect 1228 1251 1240 1252
rect 1228 1247 1232 1251
rect 1236 1247 1240 1251
rect 1429 1276 1430 1282
rect 1432 1276 1433 1282
rect 1620 1273 1621 1279
rect 1623 1273 1624 1279
rect 1790 1278 1791 1282
rect 1795 1278 1796 1282
rect 1836 1281 1837 1285
rect 1841 1281 1842 1285
rect 1746 1274 1750 1278
rect 1754 1274 1758 1278
rect 1790 1277 1796 1278
rect 1836 1280 1842 1281
rect 1873 1279 1874 1285
rect 1876 1279 1877 1285
rect 1836 1277 1842 1278
rect 1790 1274 1796 1275
rect 1746 1273 1758 1274
rect 1518 1259 1519 1265
rect 1521 1259 1522 1265
rect 1746 1270 1758 1271
rect 1790 1270 1791 1274
rect 1795 1270 1796 1274
rect 1836 1273 1837 1277
rect 1841 1273 1842 1277
rect 1746 1266 1750 1270
rect 1754 1266 1758 1270
rect 1709 1256 1710 1262
rect 1712 1256 1713 1262
rect 1746 1256 1750 1260
rect 1754 1256 1758 1260
rect 1746 1255 1758 1256
rect 1746 1252 1758 1253
rect 1746 1248 1750 1252
rect 1754 1248 1758 1252
rect 1429 1224 1430 1230
rect 1432 1224 1433 1230
rect 317 1200 318 1204
rect 322 1200 323 1204
rect 374 1203 375 1207
rect 379 1203 380 1207
rect 245 1196 249 1200
rect 253 1196 257 1200
rect 317 1199 323 1200
rect 374 1202 380 1203
rect 427 1201 428 1207
rect 430 1201 431 1207
rect 562 1204 563 1210
rect 565 1204 566 1210
rect 374 1199 380 1200
rect 317 1196 323 1197
rect 245 1195 257 1196
rect 245 1192 257 1193
rect 317 1192 318 1196
rect 322 1192 323 1196
rect 374 1195 375 1199
rect 379 1195 380 1199
rect 245 1188 249 1192
rect 253 1188 257 1192
rect 245 1178 249 1182
rect 253 1178 257 1182
rect 245 1177 257 1178
rect 245 1174 257 1175
rect 245 1170 249 1174
rect 253 1170 257 1174
rect 748 1201 749 1207
rect 751 1201 752 1207
rect 1620 1221 1621 1227
rect 1623 1221 1624 1227
rect 677 1169 678 1175
rect 680 1169 681 1175
rect 1295 1169 1296 1173
rect 1300 1169 1301 1173
rect 1341 1172 1342 1176
rect 1346 1172 1347 1176
rect 1251 1165 1255 1169
rect 1259 1165 1263 1169
rect 1295 1168 1301 1169
rect 1341 1171 1347 1172
rect 1378 1170 1379 1176
rect 1381 1170 1382 1176
rect 1341 1168 1347 1169
rect 1295 1165 1301 1166
rect 1251 1164 1263 1165
rect 1251 1161 1263 1162
rect 1295 1161 1296 1165
rect 1300 1161 1301 1165
rect 1341 1164 1342 1168
rect 1346 1164 1347 1168
rect 703 1153 704 1159
rect 706 1153 707 1159
rect 1251 1157 1255 1161
rect 1259 1157 1263 1161
rect 1251 1147 1255 1151
rect 1259 1147 1263 1151
rect 1251 1146 1263 1147
rect 1251 1143 1263 1144
rect 1251 1139 1255 1143
rect 1259 1139 1263 1143
rect 1434 1147 1435 1153
rect 1437 1147 1438 1153
rect 1460 1131 1461 1137
rect 1463 1131 1464 1137
rect 1582 1135 1583 1147
rect 1585 1135 1586 1147
rect 1769 1147 1770 1159
rect 1772 1147 1773 1159
rect 1749 1133 1750 1145
rect 1752 1133 1753 1145
rect 1872 1136 1873 1148
rect 1875 1136 1876 1148
rect 818 1112 819 1118
rect 821 1112 822 1118
rect 1730 1115 1731 1127
rect 1733 1115 1734 1127
rect 844 1096 845 1102
rect 847 1096 848 1102
rect 1479 1099 1480 1105
rect 1482 1099 1483 1105
rect 1574 1101 1575 1113
rect 1577 1101 1578 1113
rect 1605 1101 1606 1113
rect 1608 1101 1609 1113
rect 1809 1112 1810 1118
rect 1812 1112 1813 1118
rect 473 1082 474 1086
rect 478 1082 479 1086
rect 530 1085 531 1089
rect 535 1085 536 1089
rect 401 1078 405 1082
rect 409 1078 413 1082
rect 473 1081 479 1082
rect 530 1084 536 1085
rect 583 1083 584 1089
rect 586 1083 587 1089
rect 1872 1104 1873 1116
rect 1875 1104 1876 1116
rect 1905 1115 1906 1121
rect 1908 1115 1909 1121
rect 1635 1086 1636 1092
rect 1638 1086 1639 1092
rect 530 1081 536 1082
rect 473 1078 479 1079
rect 401 1077 413 1078
rect 401 1074 413 1075
rect 473 1074 474 1078
rect 478 1074 479 1078
rect 530 1077 531 1081
rect 535 1077 536 1081
rect 401 1070 405 1074
rect 409 1070 413 1074
rect 401 1060 405 1064
rect 409 1060 413 1064
rect 401 1059 413 1060
rect 401 1056 413 1057
rect 401 1052 405 1056
rect 409 1052 413 1056
rect 678 1033 679 1039
rect 681 1033 682 1039
rect 704 1017 705 1023
rect 707 1017 708 1023
rect 800 898 801 902
rect 805 898 806 902
rect 857 901 858 905
rect 862 901 863 905
rect 751 894 755 898
rect 759 894 763 898
rect 800 897 806 898
rect 857 900 863 901
rect 910 899 911 905
rect 913 899 914 905
rect 857 897 863 898
rect 800 894 806 895
rect 751 893 763 894
rect 751 890 763 891
rect 800 890 801 894
rect 805 890 806 894
rect 857 893 858 897
rect 862 893 863 897
rect 751 886 755 890
rect 759 886 763 890
rect 751 876 755 880
rect 759 876 763 880
rect 751 875 763 876
rect 751 872 763 873
rect 751 868 755 872
rect 759 868 763 872
rect 963 886 964 892
rect 966 886 967 892
rect 1124 883 1125 889
rect 1127 883 1128 889
rect 1052 869 1053 875
rect 1055 869 1056 875
rect 1308 874 1309 878
rect 1313 874 1314 878
rect 1365 877 1366 881
rect 1370 877 1371 881
rect 1213 866 1214 872
rect 1216 866 1217 872
rect 1260 870 1264 874
rect 1268 870 1272 874
rect 1308 873 1314 874
rect 1365 876 1371 877
rect 1408 875 1409 881
rect 1411 875 1412 881
rect 1365 873 1371 874
rect 1308 870 1314 871
rect 1260 869 1272 870
rect 1260 866 1272 867
rect 1308 866 1309 870
rect 1313 866 1314 870
rect 1365 869 1366 873
rect 1370 869 1371 873
rect 1260 862 1264 866
rect 1268 862 1272 866
rect 1260 852 1264 856
rect 1268 852 1272 856
rect 1260 851 1272 852
rect 1260 848 1272 849
rect 963 834 964 840
rect 966 834 967 840
rect 1260 844 1264 848
rect 1268 844 1272 848
rect 1124 831 1125 837
rect 1127 831 1128 837
rect 1717 828 1718 832
rect 1722 828 1723 832
rect 1763 831 1764 835
rect 1768 831 1769 835
rect 1673 824 1677 828
rect 1681 824 1685 828
rect 1717 827 1723 828
rect 1763 830 1769 831
rect 1800 829 1801 835
rect 1803 829 1804 835
rect 1763 827 1769 828
rect 1717 824 1723 825
rect 1673 823 1685 824
rect 1673 820 1685 821
rect 1717 820 1718 824
rect 1722 820 1723 824
rect 1763 823 1764 827
rect 1768 823 1769 827
rect 1673 816 1677 820
rect 1681 816 1685 820
rect 1673 806 1677 810
rect 1681 806 1685 810
rect 1673 805 1685 806
rect 1673 802 1685 803
rect 1673 798 1677 802
rect 1681 798 1685 802
rect 1851 816 1852 822
rect 1854 816 1855 822
rect 2111 813 2112 819
rect 2114 813 2115 819
rect 1940 799 1941 805
rect 1943 799 1944 805
rect 2281 808 2282 812
rect 2286 808 2287 812
rect 2327 811 2328 815
rect 2332 811 2333 815
rect 2237 804 2241 808
rect 2245 804 2249 808
rect 2281 807 2287 808
rect 2327 810 2333 811
rect 2364 809 2365 815
rect 2367 809 2368 815
rect 2327 807 2333 808
rect 2281 804 2287 805
rect 2237 803 2249 804
rect 2200 796 2201 802
rect 2203 796 2204 802
rect 2237 800 2249 801
rect 2281 800 2282 804
rect 2286 800 2287 804
rect 2327 803 2328 807
rect 2332 803 2333 807
rect 2237 796 2241 800
rect 2245 796 2249 800
rect 2237 786 2241 790
rect 2245 786 2249 790
rect 2237 785 2249 786
rect 2237 782 2249 783
rect 825 767 826 771
rect 830 767 831 771
rect 874 770 875 774
rect 879 770 880 774
rect 781 763 785 767
rect 789 763 793 767
rect 825 766 831 767
rect 874 769 880 770
rect 914 768 915 774
rect 917 768 918 774
rect 2237 778 2241 782
rect 2245 778 2249 782
rect 874 766 880 767
rect 825 763 831 764
rect 781 762 793 763
rect 781 759 793 760
rect 825 759 826 763
rect 830 759 831 763
rect 874 762 875 766
rect 879 762 880 766
rect 781 755 785 759
rect 789 755 793 759
rect 781 745 785 749
rect 789 745 793 749
rect 781 744 793 745
rect 781 741 793 742
rect 781 737 785 741
rect 789 737 793 741
rect 968 759 969 765
rect 971 759 972 765
rect 1116 759 1117 771
rect 1119 759 1120 771
rect 1851 764 1852 770
rect 1854 764 1855 770
rect 2111 761 2112 767
rect 2114 761 2115 767
rect 994 743 995 749
rect 997 743 998 749
rect 1108 725 1109 737
rect 1111 725 1112 737
rect 1139 725 1140 737
rect 1142 725 1143 737
rect 1013 711 1014 717
rect 1016 711 1017 717
rect 1169 710 1170 716
rect 1172 710 1173 716
rect 1717 686 1718 690
rect 1722 686 1723 690
rect 1763 689 1764 693
rect 1768 689 1769 693
rect 1673 682 1677 686
rect 1681 682 1685 686
rect 1717 685 1723 686
rect 1763 688 1769 689
rect 1800 687 1801 693
rect 1803 687 1804 693
rect 1763 685 1769 686
rect 1717 682 1723 683
rect 1673 681 1685 682
rect 1673 678 1685 679
rect 1717 678 1718 682
rect 1722 678 1723 682
rect 1763 681 1764 685
rect 1768 681 1769 685
rect 1673 674 1677 678
rect 1681 674 1685 678
rect 1673 664 1677 668
rect 1681 664 1685 668
rect 1673 663 1685 664
rect 1673 660 1685 661
rect 1673 656 1677 660
rect 1681 656 1685 660
rect 2090 681 2091 693
rect 2093 681 2094 693
rect 2073 661 2074 673
rect 2076 661 2077 673
rect 2053 647 2054 659
rect 2056 647 2057 659
rect 2191 657 2192 669
rect 2194 657 2195 669
rect 2349 669 2350 681
rect 2352 669 2353 681
rect 2329 655 2330 667
rect 2332 655 2333 667
rect 2444 658 2445 670
rect 2447 658 2448 670
rect 2573 658 2574 670
rect 2576 658 2577 670
rect 2696 664 2697 668
rect 2701 664 2702 668
rect 2742 667 2743 671
rect 2747 667 2748 671
rect 2652 660 2656 664
rect 2660 660 2664 664
rect 2696 663 2702 664
rect 2742 666 2748 667
rect 2779 665 2780 671
rect 2782 665 2783 671
rect 2742 663 2748 664
rect 2696 660 2702 661
rect 2652 659 2664 660
rect 2652 656 2664 657
rect 2696 656 2697 660
rect 2701 656 2702 660
rect 2742 659 2743 663
rect 2747 659 2748 663
rect 2652 652 2656 656
rect 2660 652 2664 656
rect 1856 628 1857 634
rect 1859 628 1860 634
rect 2034 629 2035 641
rect 2037 629 2038 641
rect 2310 637 2311 649
rect 2313 637 2314 649
rect 2183 623 2184 635
rect 2186 623 2187 635
rect 2214 623 2215 635
rect 2217 623 2218 635
rect 2385 634 2386 640
rect 2388 634 2389 640
rect 2652 642 2656 646
rect 2660 642 2664 646
rect 2652 641 2664 642
rect 2652 638 2664 639
rect 1882 612 1883 618
rect 1885 612 1886 618
rect 2444 626 2445 638
rect 2447 626 2448 638
rect 2489 625 2490 631
rect 2492 625 2493 631
rect 2573 626 2574 638
rect 2576 626 2577 638
rect 2652 634 2656 638
rect 2660 634 2664 638
rect 2244 608 2245 614
rect 2247 608 2248 614
rect 2607 625 2608 631
rect 2610 625 2611 631
rect 1905 580 1906 586
rect 1908 580 1909 586
rect 2117 522 2118 528
rect 2120 522 2121 528
<< ndcontact >>
rect 430 1278 434 1282
rect 438 1279 442 1283
rect 325 1270 329 1274
rect 382 1273 386 1277
rect 256 1260 260 1264
rect 326 1261 330 1265
rect 383 1264 387 1268
rect 256 1252 260 1256
rect 326 1245 330 1249
rect 383 1248 387 1252
rect 326 1236 330 1240
rect 383 1239 387 1243
rect 613 1250 617 1256
rect 630 1250 634 1256
rect 558 1238 562 1242
rect 566 1239 570 1243
rect 799 1247 803 1253
rect 816 1247 820 1253
rect 744 1235 748 1239
rect 752 1236 756 1240
rect 647 1221 651 1225
rect 655 1222 659 1226
rect 1480 1270 1484 1276
rect 1497 1270 1501 1276
rect 1425 1258 1429 1262
rect 1433 1259 1437 1263
rect 1671 1267 1675 1273
rect 1688 1267 1692 1273
rect 1351 1246 1355 1250
rect 1359 1247 1363 1251
rect 1273 1238 1277 1242
rect 1319 1241 1323 1245
rect 1616 1255 1620 1259
rect 1624 1256 1628 1260
rect 1514 1241 1518 1245
rect 1522 1242 1526 1246
rect 1869 1247 1873 1251
rect 1877 1248 1881 1252
rect 1705 1238 1709 1242
rect 1713 1239 1717 1243
rect 1791 1239 1795 1243
rect 1837 1242 1841 1246
rect 1047 1227 1051 1231
rect 1055 1228 1059 1232
rect 833 1218 837 1222
rect 841 1219 845 1223
rect 942 1219 946 1223
rect 999 1222 1003 1226
rect 1232 1228 1236 1232
rect 1274 1229 1278 1233
rect 1320 1232 1324 1236
rect 1480 1229 1485 1235
rect 1497 1229 1501 1235
rect 613 1209 618 1215
rect 630 1209 634 1215
rect 1232 1220 1236 1224
rect 799 1206 804 1212
rect 816 1206 820 1212
rect 873 1209 877 1213
rect 943 1210 947 1214
rect 1000 1213 1004 1217
rect 1274 1213 1278 1217
rect 1320 1216 1324 1220
rect 1671 1226 1676 1232
rect 1688 1226 1692 1232
rect 1750 1229 1754 1233
rect 1792 1230 1796 1234
rect 1838 1233 1842 1237
rect 1750 1221 1754 1225
rect 873 1201 877 1205
rect 1274 1204 1278 1208
rect 1320 1207 1324 1211
rect 1425 1206 1429 1210
rect 1433 1207 1437 1211
rect 1792 1214 1796 1218
rect 1838 1217 1842 1221
rect 1616 1203 1620 1207
rect 1624 1204 1628 1208
rect 1792 1205 1796 1209
rect 1838 1208 1842 1212
rect 558 1186 562 1190
rect 566 1187 570 1191
rect 943 1194 947 1198
rect 1000 1197 1004 1201
rect 744 1183 748 1187
rect 752 1184 756 1188
rect 943 1185 947 1189
rect 1000 1188 1004 1192
rect 423 1169 427 1173
rect 431 1170 435 1174
rect 318 1161 322 1165
rect 375 1164 379 1168
rect 249 1151 253 1155
rect 319 1152 323 1156
rect 376 1155 380 1159
rect 249 1143 253 1147
rect 319 1136 323 1140
rect 376 1139 380 1143
rect 1374 1138 1378 1142
rect 1382 1139 1386 1143
rect 319 1127 323 1131
rect 376 1130 380 1134
rect 1296 1130 1300 1134
rect 1342 1133 1346 1137
rect 681 1120 685 1126
rect 689 1120 693 1126
rect 1255 1120 1259 1124
rect 1297 1121 1301 1125
rect 1343 1124 1347 1128
rect 1255 1112 1259 1116
rect 1297 1105 1301 1109
rect 1343 1108 1347 1112
rect 681 1094 685 1100
rect 689 1094 693 1100
rect 1297 1096 1301 1100
rect 1343 1099 1347 1103
rect 1438 1098 1442 1104
rect 1446 1098 1450 1104
rect 1805 1094 1809 1098
rect 1813 1095 1817 1099
rect 1901 1097 1905 1101
rect 1909 1098 1913 1102
rect 1475 1081 1479 1085
rect 1483 1082 1487 1086
rect 1438 1072 1442 1078
rect 1446 1072 1450 1078
rect 1749 1081 1753 1090
rect 1757 1081 1761 1090
rect 1878 1080 1882 1086
rect 1886 1080 1890 1086
rect 1860 1073 1864 1079
rect 1868 1073 1872 1079
rect 822 1063 826 1069
rect 830 1063 834 1069
rect 1594 1066 1598 1072
rect 1602 1066 1606 1072
rect 1631 1068 1635 1072
rect 1639 1069 1643 1073
rect 1749 1061 1753 1070
rect 1757 1061 1761 1070
rect 579 1051 583 1055
rect 587 1052 591 1056
rect 1571 1053 1575 1059
rect 1579 1053 1583 1059
rect 474 1043 478 1047
rect 531 1046 535 1050
rect 405 1033 409 1037
rect 475 1034 479 1038
rect 532 1037 536 1041
rect 822 1037 826 1043
rect 830 1037 834 1043
rect 1594 1040 1598 1046
rect 1602 1040 1606 1046
rect 405 1025 409 1029
rect 1749 1033 1753 1042
rect 1757 1033 1761 1042
rect 475 1018 479 1022
rect 532 1021 536 1025
rect 475 1009 479 1013
rect 532 1012 536 1016
rect 682 984 686 990
rect 690 984 694 990
rect 682 958 686 964
rect 690 958 694 964
rect 1014 880 1018 886
rect 1031 880 1035 886
rect 906 867 910 871
rect 914 868 918 872
rect 959 868 963 872
rect 967 869 971 873
rect 1175 877 1179 883
rect 1192 877 1196 883
rect 801 859 805 863
rect 858 862 862 866
rect 755 849 759 853
rect 802 850 806 854
rect 859 853 863 857
rect 1120 865 1124 869
rect 1128 866 1132 870
rect 1048 851 1052 855
rect 1056 852 1060 856
rect 1209 848 1213 852
rect 1217 849 1221 853
rect 755 841 759 845
rect 802 834 806 838
rect 859 837 863 841
rect 1014 839 1019 845
rect 1031 839 1035 845
rect 1404 843 1408 847
rect 1412 844 1416 848
rect 802 825 806 829
rect 859 828 863 832
rect 1175 836 1180 842
rect 1192 836 1196 842
rect 1309 835 1313 839
rect 1366 838 1370 842
rect 959 816 963 820
rect 967 817 971 821
rect 1264 825 1268 829
rect 1310 826 1314 830
rect 1367 829 1371 833
rect 1120 813 1124 817
rect 1128 814 1132 818
rect 1264 817 1268 821
rect 1310 810 1314 814
rect 1367 813 1371 817
rect 1310 801 1314 805
rect 1367 804 1371 808
rect 1902 810 1906 816
rect 1919 810 1923 816
rect 1796 797 1800 801
rect 1804 798 1808 802
rect 1847 798 1851 802
rect 1855 799 1859 803
rect 2162 807 2166 813
rect 2179 807 2183 813
rect 1718 789 1722 793
rect 1764 792 1768 796
rect 1677 779 1681 783
rect 1719 780 1723 784
rect 1765 783 1769 787
rect 2107 795 2111 799
rect 2115 796 2119 800
rect 1936 781 1940 785
rect 1944 782 1948 786
rect 2196 778 2200 782
rect 2204 779 2208 783
rect 2360 777 2364 781
rect 2368 778 2372 782
rect 1677 771 1681 775
rect 1719 764 1723 768
rect 1765 767 1769 771
rect 1902 769 1907 775
rect 1919 769 1923 775
rect 1719 755 1723 759
rect 1765 758 1769 762
rect 2162 766 2167 772
rect 2179 766 2183 772
rect 2282 769 2286 773
rect 2328 772 2332 776
rect 2241 759 2245 763
rect 2283 760 2287 764
rect 2329 763 2333 767
rect 1847 746 1851 750
rect 1855 747 1859 751
rect 2241 751 2245 755
rect 910 736 914 740
rect 918 737 922 741
rect 2107 743 2111 747
rect 2115 744 2119 748
rect 2283 744 2287 748
rect 2329 747 2333 751
rect 826 728 830 732
rect 875 731 879 735
rect 785 718 789 722
rect 827 719 831 723
rect 876 722 880 726
rect 2283 735 2287 739
rect 2329 738 2333 742
rect 785 710 789 714
rect 972 710 976 716
rect 980 710 984 716
rect 827 703 831 707
rect 876 706 880 710
rect 827 694 831 698
rect 876 697 880 701
rect 1009 693 1013 697
rect 1017 694 1021 698
rect 1128 690 1132 696
rect 1136 690 1140 696
rect 1165 692 1169 696
rect 1173 693 1177 697
rect 972 684 976 690
rect 980 684 984 690
rect 1105 677 1109 683
rect 1113 677 1117 683
rect 1128 664 1132 670
rect 1136 664 1140 670
rect 1796 655 1800 659
rect 1804 656 1808 660
rect 1718 647 1722 651
rect 1764 650 1768 654
rect 1677 637 1681 641
rect 1719 638 1723 642
rect 1765 641 1769 645
rect 1677 629 1681 633
rect 1719 622 1723 626
rect 1765 625 1769 629
rect 1719 613 1723 617
rect 1765 616 1769 620
rect 2775 633 2779 637
rect 2783 634 2787 638
rect 2381 616 2385 620
rect 2389 617 2393 621
rect 2053 595 2057 604
rect 2061 595 2065 604
rect 2329 603 2333 612
rect 2337 603 2341 612
rect 2697 625 2701 629
rect 2743 628 2747 632
rect 2450 602 2454 608
rect 2458 602 2462 608
rect 2485 607 2489 611
rect 2493 608 2497 612
rect 2656 615 2660 619
rect 2698 616 2702 620
rect 2744 619 2748 623
rect 2432 595 2436 601
rect 2440 595 2444 601
rect 2579 602 2583 608
rect 2587 602 2591 608
rect 2603 607 2607 611
rect 2611 608 2615 612
rect 2656 607 2660 611
rect 2561 595 2565 601
rect 2569 595 2573 601
rect 2698 600 2702 604
rect 2744 603 2748 607
rect 2203 588 2207 594
rect 2211 588 2215 594
rect 2240 590 2244 594
rect 2248 591 2252 595
rect 1860 579 1864 585
rect 1868 579 1872 585
rect 2053 575 2057 584
rect 2061 575 2065 584
rect 2329 583 2333 592
rect 2337 583 2341 592
rect 2698 591 2702 595
rect 2744 594 2748 598
rect 2180 575 2184 581
rect 2188 575 2192 581
rect 1901 562 1905 566
rect 1909 563 1913 567
rect 1860 553 1864 559
rect 1868 553 1872 559
rect 2203 562 2207 568
rect 2211 562 2215 568
rect 2053 547 2057 556
rect 2061 547 2065 556
rect 2329 555 2333 564
rect 2337 555 2341 564
rect 2053 527 2057 536
rect 2061 527 2065 536
rect 2113 504 2117 508
rect 2121 505 2125 509
<< pdcontact >>
rect 325 1309 329 1313
rect 382 1312 386 1316
rect 256 1305 260 1309
rect 430 1310 434 1316
rect 438 1310 442 1316
rect 325 1301 329 1305
rect 382 1304 386 1308
rect 256 1297 260 1301
rect 256 1287 260 1291
rect 256 1279 260 1283
rect 1273 1277 1277 1281
rect 1319 1280 1323 1284
rect 1232 1273 1236 1277
rect 1351 1278 1355 1284
rect 1359 1278 1363 1284
rect 1273 1269 1277 1273
rect 1319 1272 1323 1276
rect 1232 1265 1236 1269
rect 558 1256 562 1262
rect 566 1256 570 1262
rect 744 1253 748 1259
rect 752 1253 756 1259
rect 942 1258 946 1262
rect 999 1261 1003 1265
rect 873 1254 877 1258
rect 1047 1259 1051 1265
rect 1055 1259 1059 1265
rect 647 1239 651 1245
rect 655 1239 659 1245
rect 942 1250 946 1254
rect 999 1253 1003 1257
rect 873 1246 877 1250
rect 833 1236 837 1242
rect 841 1236 845 1242
rect 873 1236 877 1240
rect 873 1228 877 1232
rect 1232 1255 1236 1259
rect 1232 1247 1236 1251
rect 1425 1276 1429 1282
rect 1433 1276 1437 1282
rect 1616 1273 1620 1279
rect 1624 1273 1628 1279
rect 1791 1278 1795 1282
rect 1837 1281 1841 1285
rect 1750 1274 1754 1278
rect 1869 1279 1873 1285
rect 1877 1279 1881 1285
rect 1514 1259 1518 1265
rect 1522 1259 1526 1265
rect 1791 1270 1795 1274
rect 1837 1273 1841 1277
rect 1750 1266 1754 1270
rect 1705 1256 1709 1262
rect 1713 1256 1717 1262
rect 1750 1256 1754 1260
rect 1750 1248 1754 1252
rect 1425 1224 1429 1230
rect 1433 1224 1437 1230
rect 318 1200 322 1204
rect 375 1203 379 1207
rect 249 1196 253 1200
rect 423 1201 427 1207
rect 431 1201 435 1207
rect 558 1204 562 1210
rect 566 1204 570 1210
rect 318 1192 322 1196
rect 375 1195 379 1199
rect 249 1188 253 1192
rect 249 1178 253 1182
rect 249 1170 253 1174
rect 744 1201 748 1207
rect 752 1201 756 1207
rect 1616 1221 1620 1227
rect 1624 1221 1628 1227
rect 673 1169 677 1175
rect 681 1169 685 1175
rect 1296 1169 1300 1173
rect 1342 1172 1346 1176
rect 1255 1165 1259 1169
rect 1374 1170 1378 1176
rect 1382 1170 1386 1176
rect 1296 1161 1300 1165
rect 1342 1164 1346 1168
rect 699 1153 703 1159
rect 707 1153 711 1159
rect 1255 1157 1259 1161
rect 1255 1147 1259 1151
rect 1255 1139 1259 1143
rect 1430 1147 1434 1153
rect 1438 1147 1442 1153
rect 1456 1131 1460 1137
rect 1464 1131 1468 1137
rect 1578 1135 1582 1147
rect 1586 1135 1590 1147
rect 1765 1147 1769 1159
rect 1773 1147 1777 1159
rect 1745 1133 1749 1145
rect 1753 1133 1757 1145
rect 1868 1136 1872 1148
rect 1876 1136 1880 1148
rect 814 1112 818 1118
rect 822 1112 826 1118
rect 1726 1115 1730 1127
rect 1734 1115 1738 1127
rect 840 1096 844 1102
rect 848 1096 852 1102
rect 1475 1099 1479 1105
rect 1483 1099 1487 1105
rect 1570 1101 1574 1113
rect 1578 1101 1582 1113
rect 1601 1101 1605 1113
rect 1609 1101 1613 1113
rect 1805 1112 1809 1118
rect 1813 1112 1817 1118
rect 474 1082 478 1086
rect 531 1085 535 1089
rect 405 1078 409 1082
rect 579 1083 583 1089
rect 587 1083 591 1089
rect 1868 1104 1872 1116
rect 1876 1104 1880 1116
rect 1901 1115 1905 1121
rect 1909 1115 1913 1121
rect 1631 1086 1635 1092
rect 1639 1086 1643 1092
rect 474 1074 478 1078
rect 531 1077 535 1081
rect 405 1070 409 1074
rect 405 1060 409 1064
rect 405 1052 409 1056
rect 674 1033 678 1039
rect 682 1033 686 1039
rect 700 1017 704 1023
rect 708 1017 712 1023
rect 801 898 805 902
rect 858 901 862 905
rect 755 894 759 898
rect 906 899 910 905
rect 914 899 918 905
rect 801 890 805 894
rect 858 893 862 897
rect 755 886 759 890
rect 755 876 759 880
rect 755 868 759 872
rect 959 886 963 892
rect 967 886 971 892
rect 1120 883 1124 889
rect 1128 883 1132 889
rect 1048 869 1052 875
rect 1056 869 1060 875
rect 1309 874 1313 878
rect 1366 877 1370 881
rect 1209 866 1213 872
rect 1217 866 1221 872
rect 1264 870 1268 874
rect 1404 875 1408 881
rect 1412 875 1416 881
rect 1309 866 1313 870
rect 1366 869 1370 873
rect 1264 862 1268 866
rect 1264 852 1268 856
rect 959 834 963 840
rect 967 834 971 840
rect 1264 844 1268 848
rect 1120 831 1124 837
rect 1128 831 1132 837
rect 1718 828 1722 832
rect 1764 831 1768 835
rect 1677 824 1681 828
rect 1796 829 1800 835
rect 1804 829 1808 835
rect 1718 820 1722 824
rect 1764 823 1768 827
rect 1677 816 1681 820
rect 1677 806 1681 810
rect 1677 798 1681 802
rect 1847 816 1851 822
rect 1855 816 1859 822
rect 2107 813 2111 819
rect 2115 813 2119 819
rect 1936 799 1940 805
rect 1944 799 1948 805
rect 2282 808 2286 812
rect 2328 811 2332 815
rect 2241 804 2245 808
rect 2360 809 2364 815
rect 2368 809 2372 815
rect 2196 796 2200 802
rect 2204 796 2208 802
rect 2282 800 2286 804
rect 2328 803 2332 807
rect 2241 796 2245 800
rect 2241 786 2245 790
rect 826 767 830 771
rect 875 770 879 774
rect 785 763 789 767
rect 910 768 914 774
rect 918 768 922 774
rect 2241 778 2245 782
rect 826 759 830 763
rect 875 762 879 766
rect 785 755 789 759
rect 785 745 789 749
rect 785 737 789 741
rect 964 759 968 765
rect 972 759 976 765
rect 1112 759 1116 771
rect 1120 759 1124 771
rect 1847 764 1851 770
rect 1855 764 1859 770
rect 2107 761 2111 767
rect 2115 761 2119 767
rect 990 743 994 749
rect 998 743 1002 749
rect 1104 725 1108 737
rect 1112 725 1116 737
rect 1135 725 1139 737
rect 1143 725 1147 737
rect 1009 711 1013 717
rect 1017 711 1021 717
rect 1165 710 1169 716
rect 1173 710 1177 716
rect 1718 686 1722 690
rect 1764 689 1768 693
rect 1677 682 1681 686
rect 1796 687 1800 693
rect 1804 687 1808 693
rect 1718 678 1722 682
rect 1764 681 1768 685
rect 1677 674 1681 678
rect 1677 664 1681 668
rect 1677 656 1681 660
rect 2086 681 2090 693
rect 2094 681 2098 693
rect 2069 661 2073 673
rect 2077 661 2081 673
rect 2049 647 2053 659
rect 2057 647 2061 659
rect 2187 657 2191 669
rect 2195 657 2199 669
rect 2345 669 2349 681
rect 2353 669 2357 681
rect 2325 655 2329 667
rect 2333 655 2337 667
rect 2440 658 2444 670
rect 2448 658 2452 670
rect 2569 658 2573 670
rect 2577 658 2581 670
rect 2697 664 2701 668
rect 2743 667 2747 671
rect 2656 660 2660 664
rect 2775 665 2779 671
rect 2783 665 2787 671
rect 2697 656 2701 660
rect 2743 659 2747 663
rect 2656 652 2660 656
rect 1852 628 1856 634
rect 1860 628 1864 634
rect 2030 629 2034 641
rect 2038 629 2042 641
rect 2306 637 2310 649
rect 2314 637 2318 649
rect 2179 623 2183 635
rect 2187 623 2191 635
rect 2210 623 2214 635
rect 2218 623 2222 635
rect 2381 634 2385 640
rect 2389 634 2393 640
rect 2656 642 2660 646
rect 1878 612 1882 618
rect 1886 612 1890 618
rect 2440 626 2444 638
rect 2448 626 2452 638
rect 2485 625 2489 631
rect 2493 625 2497 631
rect 2569 626 2573 638
rect 2577 626 2581 638
rect 2656 634 2660 638
rect 2240 608 2244 614
rect 2248 608 2252 614
rect 2603 625 2607 631
rect 2611 625 2615 631
rect 1901 580 1905 586
rect 1909 580 1913 586
rect 2113 522 2117 528
rect 2121 522 2125 528
<< polysilicon >>
rect 435 1316 437 1319
rect 375 1309 381 1311
rect 387 1309 395 1311
rect 318 1306 324 1308
rect 330 1306 338 1308
rect 245 1302 252 1304
rect 264 1302 271 1304
rect 245 1284 252 1286
rect 264 1284 271 1286
rect 435 1282 437 1310
rect 1356 1284 1358 1287
rect 1874 1285 1876 1288
rect 435 1276 437 1279
rect 1312 1277 1318 1279
rect 1324 1277 1332 1279
rect 1430 1282 1432 1285
rect 1266 1274 1272 1276
rect 1278 1274 1286 1276
rect 374 1269 382 1271
rect 388 1269 394 1271
rect 1221 1270 1228 1272
rect 1240 1270 1247 1272
rect 317 1266 325 1268
rect 331 1266 337 1268
rect 1052 1265 1054 1268
rect 563 1262 565 1265
rect 245 1257 257 1259
rect 260 1257 271 1259
rect 749 1259 751 1262
rect 622 1256 624 1259
rect 374 1244 382 1246
rect 388 1244 394 1246
rect 317 1241 325 1243
rect 331 1241 337 1243
rect 563 1242 565 1256
rect 808 1253 810 1256
rect 992 1258 998 1260
rect 1004 1258 1012 1260
rect 935 1255 941 1257
rect 947 1255 955 1257
rect 622 1241 624 1250
rect 652 1245 654 1248
rect 749 1239 751 1253
rect 862 1251 869 1253
rect 881 1251 888 1253
rect 563 1236 565 1239
rect 652 1225 654 1239
rect 808 1238 810 1247
rect 838 1242 840 1245
rect 749 1233 751 1236
rect 838 1222 840 1236
rect 862 1233 869 1235
rect 881 1233 888 1235
rect 1052 1231 1054 1259
rect 1221 1252 1228 1254
rect 1240 1252 1247 1254
rect 1356 1250 1358 1278
rect 1621 1279 1623 1282
rect 1489 1276 1491 1279
rect 1430 1262 1432 1276
rect 1680 1273 1682 1276
rect 1830 1278 1836 1280
rect 1842 1278 1850 1280
rect 1784 1275 1790 1277
rect 1796 1275 1804 1277
rect 1489 1261 1491 1270
rect 1519 1265 1521 1268
rect 1621 1259 1623 1273
rect 1739 1271 1746 1273
rect 1758 1271 1765 1273
rect 1430 1256 1432 1259
rect 1356 1244 1358 1247
rect 1519 1245 1521 1259
rect 1680 1258 1682 1267
rect 1710 1262 1712 1265
rect 1621 1253 1623 1256
rect 1710 1242 1712 1256
rect 1739 1253 1746 1255
rect 1758 1253 1765 1255
rect 1874 1251 1876 1279
rect 1519 1239 1521 1242
rect 1311 1237 1319 1239
rect 1325 1237 1331 1239
rect 1874 1245 1876 1248
rect 1265 1234 1273 1236
rect 1279 1234 1285 1236
rect 652 1219 654 1222
rect 1052 1225 1054 1228
rect 1489 1235 1491 1238
rect 1710 1236 1712 1239
rect 1430 1230 1432 1233
rect 1221 1225 1233 1227
rect 1236 1225 1247 1227
rect 1680 1232 1682 1235
rect 1829 1238 1837 1240
rect 1843 1238 1849 1240
rect 1783 1235 1791 1237
rect 1797 1235 1803 1237
rect 622 1215 624 1218
rect 838 1216 840 1219
rect 563 1210 565 1213
rect 428 1207 430 1210
rect 368 1200 374 1202
rect 380 1200 388 1202
rect 808 1212 810 1215
rect 991 1218 999 1220
rect 1005 1218 1011 1220
rect 934 1215 942 1217
rect 948 1215 954 1217
rect 311 1197 317 1199
rect 323 1197 331 1199
rect 238 1193 245 1195
rect 257 1193 264 1195
rect 238 1175 245 1177
rect 257 1175 264 1177
rect 428 1173 430 1201
rect 563 1197 565 1204
rect 622 1200 624 1209
rect 749 1207 751 1210
rect 1430 1217 1432 1224
rect 1489 1220 1491 1229
rect 1621 1227 1623 1230
rect 1739 1226 1751 1228
rect 1754 1226 1765 1228
rect 1311 1212 1319 1214
rect 1325 1212 1331 1214
rect 1429 1213 1432 1217
rect 1621 1214 1623 1221
rect 1680 1217 1682 1226
rect 1265 1209 1273 1211
rect 1279 1209 1285 1211
rect 862 1206 874 1208
rect 877 1206 888 1208
rect 562 1193 565 1197
rect 749 1194 751 1201
rect 808 1197 810 1206
rect 1430 1210 1432 1213
rect 1620 1210 1623 1214
rect 1621 1207 1623 1210
rect 1829 1213 1837 1215
rect 1843 1213 1849 1215
rect 1783 1210 1791 1212
rect 1797 1210 1803 1212
rect 1430 1204 1432 1207
rect 1621 1201 1623 1204
rect 563 1190 565 1193
rect 748 1190 751 1194
rect 749 1187 751 1190
rect 991 1193 999 1195
rect 1005 1193 1011 1195
rect 934 1190 942 1192
rect 948 1190 954 1192
rect 563 1184 565 1187
rect 749 1181 751 1184
rect 678 1175 680 1178
rect 1379 1176 1381 1179
rect 428 1167 430 1170
rect 678 1162 680 1169
rect 367 1160 375 1162
rect 381 1160 387 1162
rect 704 1159 706 1166
rect 1335 1169 1341 1171
rect 1347 1169 1355 1171
rect 1289 1166 1295 1168
rect 1301 1166 1309 1168
rect 1244 1162 1251 1164
rect 1263 1162 1270 1164
rect 310 1157 318 1159
rect 324 1157 330 1159
rect 704 1150 706 1153
rect 238 1148 250 1150
rect 253 1148 264 1150
rect 1244 1144 1251 1146
rect 1263 1144 1270 1146
rect 1379 1142 1381 1170
rect 1770 1159 1772 1166
rect 1435 1153 1437 1156
rect 1583 1147 1585 1154
rect 1435 1140 1437 1147
rect 367 1135 375 1137
rect 381 1135 387 1137
rect 310 1132 318 1134
rect 324 1132 330 1134
rect 686 1126 688 1133
rect 1379 1136 1381 1139
rect 1461 1137 1463 1144
rect 1750 1145 1752 1152
rect 1873 1148 1875 1155
rect 1583 1132 1585 1135
rect 1334 1129 1342 1131
rect 1348 1129 1354 1131
rect 1461 1128 1463 1131
rect 1288 1126 1296 1128
rect 1302 1126 1308 1128
rect 686 1117 688 1120
rect 819 1118 821 1121
rect 1731 1127 1733 1134
rect 1770 1144 1772 1147
rect 1873 1133 1875 1136
rect 1750 1130 1752 1133
rect 1244 1117 1256 1119
rect 1259 1117 1270 1119
rect 1575 1113 1577 1120
rect 1606 1113 1608 1116
rect 1810 1118 1812 1121
rect 819 1105 821 1112
rect 686 1100 688 1103
rect 845 1102 847 1109
rect 1334 1104 1342 1106
rect 1348 1104 1354 1106
rect 1443 1104 1445 1111
rect 1480 1105 1482 1108
rect 1288 1101 1296 1103
rect 1302 1101 1308 1103
rect 1731 1112 1733 1115
rect 1873 1116 1875 1123
rect 1906 1121 1908 1124
rect 584 1089 586 1092
rect 524 1082 530 1084
rect 536 1082 544 1084
rect 686 1087 688 1094
rect 845 1093 847 1096
rect 1443 1095 1445 1098
rect 1480 1085 1482 1099
rect 1575 1098 1577 1101
rect 1606 1094 1608 1101
rect 1810 1098 1812 1112
rect 1873 1101 1875 1104
rect 1906 1101 1908 1115
rect 1636 1092 1638 1095
rect 1754 1090 1756 1097
rect 1906 1095 1908 1098
rect 1810 1092 1812 1095
rect 467 1079 473 1081
rect 479 1079 487 1081
rect 394 1075 401 1077
rect 413 1075 420 1077
rect 394 1057 401 1059
rect 413 1057 420 1059
rect 584 1055 586 1083
rect 1443 1078 1445 1081
rect 1480 1079 1482 1082
rect 827 1069 829 1076
rect 1599 1072 1601 1079
rect 1636 1072 1638 1086
rect 1883 1086 1885 1089
rect 1754 1078 1756 1081
rect 1865 1079 1867 1086
rect 1883 1073 1885 1080
rect 1443 1065 1445 1072
rect 1754 1070 1756 1073
rect 1865 1070 1867 1073
rect 1636 1066 1638 1069
rect 1599 1063 1601 1066
rect 827 1060 829 1063
rect 1576 1059 1578 1062
rect 1754 1054 1756 1061
rect 584 1049 586 1052
rect 1576 1046 1578 1053
rect 1599 1046 1601 1049
rect 523 1042 531 1044
rect 537 1042 543 1044
rect 827 1043 829 1046
rect 466 1039 474 1041
rect 480 1039 486 1041
rect 679 1039 681 1042
rect 1754 1042 1756 1049
rect 394 1030 406 1032
rect 409 1030 420 1032
rect 679 1026 681 1033
rect 827 1030 829 1037
rect 1599 1033 1601 1040
rect 1754 1030 1756 1033
rect 705 1023 707 1030
rect 523 1017 531 1019
rect 537 1017 543 1019
rect 466 1014 474 1016
rect 480 1014 486 1016
rect 705 1014 707 1017
rect 687 990 689 997
rect 687 981 689 984
rect 687 964 689 967
rect 687 951 689 958
rect 911 905 913 908
rect 851 898 857 900
rect 863 898 871 900
rect 794 895 800 897
rect 806 895 814 897
rect 744 891 751 893
rect 763 891 770 893
rect 744 873 751 875
rect 763 873 770 875
rect 911 871 913 899
rect 964 892 966 895
rect 1125 889 1127 892
rect 1023 886 1025 889
rect 964 872 966 886
rect 1184 883 1186 886
rect 1023 871 1025 880
rect 1053 875 1055 878
rect 1125 869 1127 883
rect 1409 881 1411 884
rect 911 865 913 868
rect 964 866 966 869
rect 850 858 858 860
rect 864 858 870 860
rect 793 855 801 857
rect 807 855 813 857
rect 1053 855 1055 869
rect 1184 868 1186 877
rect 1214 872 1216 875
rect 1359 874 1365 876
rect 1371 874 1379 876
rect 1302 871 1308 873
rect 1314 871 1322 873
rect 1253 867 1260 869
rect 1272 867 1279 869
rect 1125 863 1127 866
rect 1214 852 1216 866
rect 1053 849 1055 852
rect 1253 849 1260 851
rect 1272 849 1279 851
rect 744 846 756 848
rect 759 846 770 848
rect 1023 845 1025 848
rect 1214 846 1216 849
rect 964 840 966 843
rect 850 833 858 835
rect 864 833 870 835
rect 1184 842 1186 845
rect 1409 847 1411 875
rect 793 830 801 832
rect 807 830 813 832
rect 964 827 966 834
rect 1023 830 1025 839
rect 1125 837 1127 840
rect 963 823 966 827
rect 1125 824 1127 831
rect 1184 827 1186 836
rect 1409 841 1411 844
rect 1358 834 1366 836
rect 1372 834 1378 836
rect 1801 835 1803 838
rect 1301 831 1309 833
rect 1315 831 1321 833
rect 964 820 966 823
rect 1124 820 1127 824
rect 1253 822 1265 824
rect 1268 822 1279 824
rect 1757 828 1763 830
rect 1769 828 1777 830
rect 1711 825 1717 827
rect 1723 825 1731 827
rect 1666 821 1673 823
rect 1685 821 1692 823
rect 1125 817 1127 820
rect 964 814 966 817
rect 1125 811 1127 814
rect 1358 809 1366 811
rect 1372 809 1378 811
rect 1301 806 1309 808
rect 1315 806 1321 808
rect 1666 803 1673 805
rect 1685 803 1692 805
rect 1801 801 1803 829
rect 1852 822 1854 825
rect 2112 819 2114 822
rect 1911 816 1913 819
rect 1852 802 1854 816
rect 2171 813 2173 816
rect 2365 815 2367 818
rect 1911 801 1913 810
rect 1941 805 1943 808
rect 2112 799 2114 813
rect 1801 795 1803 798
rect 1852 796 1854 799
rect 1756 788 1764 790
rect 1770 788 1776 790
rect 1710 785 1718 787
rect 1724 785 1730 787
rect 1941 785 1943 799
rect 2171 798 2173 807
rect 2201 802 2203 805
rect 2321 808 2327 810
rect 2333 808 2341 810
rect 2275 805 2281 807
rect 2287 805 2295 807
rect 2230 801 2237 803
rect 2249 801 2256 803
rect 2112 793 2114 796
rect 2201 782 2203 796
rect 2230 783 2237 785
rect 2249 783 2256 785
rect 1941 779 1943 782
rect 915 774 917 777
rect 868 767 874 769
rect 880 767 888 769
rect 1117 771 1119 778
rect 1666 776 1678 778
rect 1681 776 1692 778
rect 1911 775 1913 778
rect 2201 776 2203 779
rect 2365 781 2367 809
rect 819 764 825 766
rect 831 764 839 766
rect 774 760 781 762
rect 793 760 800 762
rect 774 742 781 744
rect 793 742 800 744
rect 915 740 917 768
rect 969 765 971 768
rect 1852 770 1854 773
rect 1756 763 1764 765
rect 1770 763 1776 765
rect 2171 772 2173 775
rect 1710 760 1718 762
rect 1724 760 1730 762
rect 969 752 971 759
rect 1117 756 1119 759
rect 995 749 997 756
rect 1852 757 1854 764
rect 1911 760 1913 769
rect 2112 767 2114 770
rect 2365 775 2367 778
rect 1851 753 1854 757
rect 2112 754 2114 761
rect 2171 757 2173 766
rect 2320 768 2328 770
rect 2334 768 2340 770
rect 2274 765 2282 767
rect 2288 765 2294 767
rect 2230 756 2242 758
rect 2245 756 2256 758
rect 1852 750 1854 753
rect 2111 750 2114 754
rect 2112 747 2114 750
rect 1852 744 1854 747
rect 995 740 997 743
rect 1109 737 1111 744
rect 2112 741 2114 744
rect 1140 737 1142 740
rect 2320 743 2328 745
rect 2334 743 2340 745
rect 2274 740 2282 742
rect 2288 740 2294 742
rect 915 734 917 737
rect 867 727 875 729
rect 881 727 887 729
rect 818 724 826 726
rect 832 724 838 726
rect 774 715 786 717
rect 789 715 800 717
rect 977 716 979 723
rect 1109 722 1111 725
rect 1014 717 1016 720
rect 1140 718 1142 725
rect 1170 716 1172 719
rect 977 707 979 710
rect 867 702 875 704
rect 881 702 887 704
rect 818 699 826 701
rect 832 699 838 701
rect 1014 697 1016 711
rect 1133 696 1135 703
rect 1170 696 1172 710
rect 977 690 979 693
rect 1014 691 1016 694
rect 1801 693 1803 696
rect 2091 693 2093 700
rect 1170 690 1172 693
rect 1133 687 1135 690
rect 977 677 979 684
rect 1110 683 1112 686
rect 1757 686 1763 688
rect 1769 686 1777 688
rect 1711 683 1717 685
rect 1723 683 1731 685
rect 1666 679 1673 681
rect 1685 679 1692 681
rect 1110 670 1112 677
rect 1133 670 1135 673
rect 1133 657 1135 664
rect 1666 661 1673 663
rect 1685 661 1692 663
rect 1801 659 1803 687
rect 2350 681 2352 688
rect 2074 673 2076 680
rect 2091 678 2093 681
rect 2054 659 2056 666
rect 2192 669 2194 676
rect 1801 653 1803 656
rect 1756 646 1764 648
rect 1770 646 1776 648
rect 1710 643 1718 645
rect 1724 643 1730 645
rect 2035 641 2037 648
rect 2074 658 2076 661
rect 2330 667 2332 674
rect 2445 670 2447 677
rect 2574 670 2576 677
rect 2780 671 2782 674
rect 2192 654 2194 657
rect 2311 649 2313 656
rect 2350 666 2352 669
rect 2736 664 2742 666
rect 2748 664 2756 666
rect 2690 661 2696 663
rect 2702 661 2710 663
rect 2445 655 2447 658
rect 2574 655 2576 658
rect 2645 657 2652 659
rect 2664 657 2671 659
rect 2330 652 2332 655
rect 2054 644 2056 647
rect 1666 634 1678 636
rect 1681 634 1692 636
rect 1857 634 1859 637
rect 2184 635 2186 642
rect 2215 635 2217 638
rect 2386 640 2388 643
rect 1756 621 1764 623
rect 1770 621 1776 623
rect 1857 621 1859 628
rect 2035 626 2037 629
rect 1710 618 1718 620
rect 1724 618 1730 620
rect 1883 618 1885 625
rect 2311 634 2313 637
rect 2445 638 2447 645
rect 2574 638 2576 645
rect 2645 639 2652 641
rect 2664 639 2671 641
rect 2184 620 2186 623
rect 2215 616 2217 623
rect 2386 620 2388 634
rect 2490 631 2492 634
rect 2445 623 2447 626
rect 2780 637 2782 665
rect 2608 631 2610 634
rect 2245 614 2247 617
rect 1883 609 1885 612
rect 2058 604 2060 611
rect 2334 612 2336 619
rect 2386 614 2388 617
rect 2058 592 2060 595
rect 2208 594 2210 601
rect 2245 594 2247 608
rect 2490 611 2492 625
rect 2574 623 2576 626
rect 2780 631 2782 634
rect 2455 608 2457 611
rect 2334 600 2336 603
rect 2437 601 2439 608
rect 2608 611 2610 625
rect 2735 624 2743 626
rect 2749 624 2755 626
rect 2689 621 2697 623
rect 2703 621 2709 623
rect 2645 612 2657 614
rect 2660 612 2671 614
rect 2584 608 2586 611
rect 2490 605 2492 608
rect 2455 595 2457 602
rect 2566 601 2568 608
rect 2608 605 2610 608
rect 2584 595 2586 602
rect 2735 599 2743 601
rect 2749 599 2755 601
rect 2689 596 2697 598
rect 2703 596 2709 598
rect 1865 585 1867 592
rect 1906 586 1908 589
rect 2334 592 2336 595
rect 2437 592 2439 595
rect 2566 592 2568 595
rect 2245 588 2247 591
rect 2058 584 2060 587
rect 2208 585 2210 588
rect 1865 576 1867 579
rect 1906 566 1908 580
rect 2185 581 2187 584
rect 2334 576 2336 583
rect 2058 568 2060 575
rect 2185 568 2187 575
rect 2208 568 2210 571
rect 1865 559 1867 562
rect 1906 560 1908 563
rect 2058 556 2060 563
rect 2334 564 2336 571
rect 1865 546 1867 553
rect 2208 555 2210 562
rect 2334 552 2336 555
rect 2058 544 2060 547
rect 2058 536 2060 539
rect 2118 528 2120 531
rect 2058 520 2060 527
rect 2118 508 2120 522
rect 2118 502 2120 505
<< polycontact >>
rect 245 1304 249 1308
rect 314 1305 318 1309
rect 371 1308 375 1312
rect 245 1286 249 1290
rect 431 1286 435 1290
rect 313 1265 317 1269
rect 370 1268 374 1272
rect 1221 1272 1225 1276
rect 1262 1273 1266 1277
rect 1308 1276 1312 1280
rect 245 1259 249 1263
rect 313 1240 317 1244
rect 370 1243 374 1247
rect 559 1245 563 1249
rect 862 1253 866 1257
rect 931 1254 935 1258
rect 988 1257 992 1261
rect 618 1241 622 1246
rect 745 1242 749 1246
rect 648 1228 652 1232
rect 804 1238 808 1243
rect 834 1225 838 1229
rect 862 1235 866 1239
rect 1048 1235 1052 1239
rect 1221 1254 1225 1258
rect 1352 1254 1356 1258
rect 1426 1265 1430 1269
rect 1739 1273 1743 1277
rect 1780 1274 1784 1278
rect 1826 1277 1830 1281
rect 1485 1261 1489 1266
rect 1617 1262 1621 1266
rect 1515 1248 1519 1252
rect 1676 1258 1680 1263
rect 1706 1245 1710 1249
rect 1739 1255 1743 1259
rect 1870 1255 1874 1259
rect 1261 1233 1265 1237
rect 1307 1236 1311 1240
rect 1221 1227 1225 1231
rect 1779 1234 1783 1238
rect 1825 1237 1829 1241
rect 238 1195 242 1199
rect 307 1196 311 1200
rect 364 1199 368 1203
rect 930 1214 934 1218
rect 987 1217 991 1221
rect 238 1177 242 1181
rect 424 1177 428 1181
rect 618 1200 622 1204
rect 862 1208 866 1212
rect 1485 1220 1489 1224
rect 1739 1228 1743 1232
rect 1261 1208 1265 1212
rect 1307 1211 1311 1215
rect 1425 1213 1429 1217
rect 1676 1217 1680 1221
rect 558 1193 562 1197
rect 804 1197 808 1201
rect 1616 1210 1620 1214
rect 1779 1209 1783 1213
rect 1825 1212 1829 1216
rect 744 1190 748 1194
rect 930 1189 934 1193
rect 987 1192 991 1196
rect 306 1156 310 1160
rect 363 1159 367 1163
rect 674 1162 678 1166
rect 700 1162 704 1166
rect 1244 1164 1248 1168
rect 1285 1165 1289 1169
rect 1331 1168 1335 1172
rect 238 1150 242 1154
rect 1244 1146 1248 1150
rect 1375 1146 1379 1150
rect 1766 1162 1770 1166
rect 1579 1150 1583 1154
rect 1746 1148 1750 1152
rect 306 1131 310 1135
rect 363 1134 367 1138
rect 1431 1140 1435 1144
rect 1457 1140 1461 1144
rect 682 1129 686 1133
rect 1284 1125 1288 1129
rect 1330 1128 1334 1132
rect 1869 1151 1873 1155
rect 1727 1130 1731 1134
rect 1244 1119 1248 1123
rect 1571 1116 1575 1120
rect 1869 1119 1873 1123
rect 815 1105 819 1109
rect 841 1105 845 1109
rect 1284 1100 1288 1104
rect 1330 1103 1334 1107
rect 1439 1107 1443 1111
rect 1806 1101 1810 1105
rect 394 1077 398 1081
rect 463 1078 467 1082
rect 520 1081 524 1085
rect 682 1087 686 1091
rect 1476 1088 1480 1092
rect 1602 1094 1606 1098
rect 1902 1104 1906 1108
rect 1750 1093 1754 1097
rect 394 1059 398 1063
rect 580 1059 584 1063
rect 823 1072 827 1076
rect 1595 1075 1599 1079
rect 1632 1075 1636 1079
rect 1861 1082 1865 1086
rect 1879 1073 1883 1077
rect 1439 1065 1443 1069
rect 1750 1054 1754 1058
rect 1572 1046 1576 1050
rect 462 1038 466 1042
rect 519 1041 523 1045
rect 394 1032 398 1036
rect 1750 1045 1754 1049
rect 675 1026 679 1030
rect 823 1030 827 1034
rect 1595 1033 1599 1037
rect 701 1026 705 1030
rect 462 1013 466 1017
rect 519 1016 523 1020
rect 683 993 687 997
rect 683 951 687 955
rect 744 893 748 897
rect 790 894 794 898
rect 847 897 851 901
rect 744 875 748 879
rect 907 875 911 879
rect 960 875 964 879
rect 1019 871 1023 876
rect 1121 872 1125 876
rect 789 854 793 858
rect 846 857 850 861
rect 1049 858 1053 862
rect 744 848 748 852
rect 1180 868 1184 873
rect 1253 869 1257 873
rect 1298 870 1302 874
rect 1355 873 1359 877
rect 1210 855 1214 859
rect 1253 851 1257 855
rect 1405 851 1409 855
rect 789 829 793 833
rect 846 832 850 836
rect 1019 830 1023 834
rect 959 823 963 827
rect 1180 827 1184 831
rect 1297 830 1301 834
rect 1354 833 1358 837
rect 1120 820 1124 824
rect 1253 824 1257 828
rect 1666 823 1670 827
rect 1707 824 1711 828
rect 1753 827 1757 831
rect 1297 805 1301 809
rect 1354 808 1358 812
rect 1666 805 1670 809
rect 1797 805 1801 809
rect 1848 805 1852 809
rect 1907 801 1911 806
rect 2108 802 2112 806
rect 1706 784 1710 788
rect 1752 787 1756 791
rect 1937 788 1941 792
rect 1666 778 1670 782
rect 2167 798 2171 803
rect 2230 803 2234 807
rect 2271 804 2275 808
rect 2317 807 2321 811
rect 2197 785 2201 789
rect 2230 785 2234 789
rect 2361 785 2365 789
rect 1113 774 1117 778
rect 774 762 778 766
rect 815 763 819 767
rect 864 766 868 770
rect 774 744 778 748
rect 911 744 915 748
rect 1706 759 1710 763
rect 1752 762 1756 766
rect 965 752 969 756
rect 991 752 995 756
rect 1907 760 1911 764
rect 1847 753 1851 757
rect 2167 757 2171 761
rect 2270 764 2274 768
rect 2316 767 2320 771
rect 2230 758 2234 762
rect 2107 750 2111 754
rect 1105 740 1109 744
rect 2270 739 2274 743
rect 2316 742 2320 746
rect 814 723 818 727
rect 863 726 867 730
rect 774 717 778 721
rect 973 719 977 723
rect 1136 718 1140 722
rect 814 698 818 702
rect 863 701 867 705
rect 1010 700 1014 704
rect 1129 699 1133 703
rect 1166 699 1170 703
rect 2087 696 2091 700
rect 973 677 977 681
rect 1666 681 1670 685
rect 1707 682 1711 686
rect 1753 685 1757 689
rect 1106 670 1110 674
rect 1129 657 1133 661
rect 1666 663 1670 667
rect 1797 663 1801 667
rect 2346 684 2350 688
rect 2070 676 2074 680
rect 2050 662 2054 666
rect 2188 672 2192 676
rect 2326 670 2330 674
rect 1706 642 1710 646
rect 1752 645 1756 649
rect 1666 636 1670 640
rect 2031 644 2035 648
rect 2441 673 2445 677
rect 2570 673 2574 677
rect 2307 652 2311 656
rect 2645 659 2649 663
rect 2686 660 2690 664
rect 2732 663 2736 667
rect 2180 638 2184 642
rect 2441 641 2445 645
rect 1706 617 1710 621
rect 1752 620 1756 624
rect 1853 621 1857 625
rect 1879 621 1883 625
rect 2570 641 2574 645
rect 2645 641 2649 645
rect 2776 641 2780 645
rect 2382 623 2386 627
rect 2211 616 2215 620
rect 2330 615 2334 619
rect 2054 607 2058 611
rect 2486 614 2490 618
rect 2204 597 2208 601
rect 2241 597 2245 601
rect 2604 614 2608 618
rect 2433 604 2437 608
rect 2685 620 2689 624
rect 2731 623 2735 627
rect 2645 614 2649 618
rect 2562 604 2566 608
rect 2451 595 2455 599
rect 2580 595 2584 599
rect 2685 595 2689 599
rect 2731 598 2735 602
rect 1861 588 1865 592
rect 1902 569 1906 573
rect 2330 576 2334 580
rect 2054 568 2058 572
rect 2181 568 2185 572
rect 2054 559 2058 563
rect 2330 567 2334 571
rect 1861 546 1865 550
rect 2204 555 2208 559
rect 2054 520 2058 524
rect 2114 511 2118 515
<< metal1 >>
rect 342 1324 448 1327
rect 273 1323 448 1324
rect 273 1320 346 1323
rect 367 1322 448 1323
rect 367 1320 401 1322
rect 273 1319 277 1320
rect 240 1315 277 1319
rect 310 1318 346 1320
rect 256 1309 260 1315
rect 325 1313 329 1318
rect 382 1316 386 1320
rect 430 1316 434 1322
rect 351 1308 371 1312
rect 256 1291 260 1297
rect 256 1269 260 1279
rect 325 1282 329 1301
rect 351 1282 355 1308
rect 325 1278 355 1282
rect 325 1274 329 1278
rect 256 1265 313 1269
rect 256 1264 260 1265
rect 240 1248 274 1252
rect 270 1232 274 1248
rect 326 1249 330 1261
rect 351 1247 355 1278
rect 382 1285 386 1304
rect 438 1290 442 1310
rect 1410 1296 1484 1301
rect 1290 1292 1369 1295
rect 1249 1291 1369 1292
rect 417 1286 431 1290
rect 438 1286 518 1290
rect 1249 1288 1294 1291
rect 1304 1290 1369 1291
rect 1304 1288 1338 1290
rect 1249 1287 1253 1288
rect 417 1285 421 1286
rect 382 1281 421 1285
rect 438 1283 442 1286
rect 382 1277 386 1281
rect 430 1268 434 1278
rect 383 1252 387 1264
rect 423 1264 434 1268
rect 351 1243 370 1247
rect 326 1232 330 1236
rect 383 1235 387 1239
rect 423 1235 427 1264
rect 369 1232 427 1235
rect 270 1231 427 1232
rect 270 1228 373 1231
rect 335 1215 441 1218
rect 266 1214 441 1215
rect 266 1211 339 1214
rect 360 1213 441 1214
rect 360 1211 394 1213
rect 266 1210 270 1211
rect 233 1206 270 1210
rect 303 1209 339 1211
rect 249 1200 253 1206
rect 318 1204 322 1209
rect 375 1207 379 1211
rect 423 1207 427 1213
rect 344 1199 364 1203
rect 249 1182 253 1188
rect 249 1160 253 1170
rect 318 1173 322 1192
rect 344 1173 348 1199
rect 318 1169 348 1173
rect 318 1165 322 1169
rect 249 1156 306 1160
rect 249 1155 253 1156
rect 233 1139 267 1143
rect 263 1123 267 1139
rect 319 1140 323 1152
rect 344 1138 348 1169
rect 375 1176 379 1195
rect 431 1181 435 1201
rect 410 1177 424 1181
rect 431 1177 438 1181
rect 410 1176 414 1177
rect 375 1172 414 1176
rect 431 1174 435 1177
rect 375 1168 379 1172
rect 423 1159 427 1169
rect 376 1143 380 1155
rect 416 1155 427 1159
rect 344 1134 363 1138
rect 319 1123 323 1127
rect 376 1126 380 1130
rect 416 1126 420 1155
rect 470 1145 474 1286
rect 514 1249 518 1286
rect 1216 1283 1253 1287
rect 1258 1286 1294 1288
rect 543 1276 617 1281
rect 543 1249 547 1276
rect 552 1267 576 1271
rect 558 1262 562 1267
rect 613 1256 617 1276
rect 729 1273 803 1278
rect 1232 1277 1236 1283
rect 1273 1281 1277 1286
rect 1319 1284 1323 1288
rect 1351 1284 1355 1290
rect 959 1273 1065 1276
rect 641 1250 665 1254
rect 514 1245 559 1249
rect 558 1235 562 1238
rect 552 1231 576 1235
rect 630 1232 634 1250
rect 647 1245 651 1250
rect 729 1246 733 1273
rect 738 1264 762 1268
rect 744 1259 748 1264
rect 799 1253 803 1273
rect 890 1272 1065 1273
rect 1299 1276 1308 1280
rect 890 1269 963 1272
rect 984 1271 1065 1272
rect 984 1269 1018 1271
rect 890 1268 894 1269
rect 857 1264 894 1268
rect 927 1267 963 1269
rect 873 1258 877 1264
rect 942 1262 946 1267
rect 999 1265 1003 1269
rect 1047 1265 1051 1271
rect 854 1253 862 1257
rect 968 1257 988 1261
rect 827 1247 851 1251
rect 655 1233 659 1239
rect 708 1242 745 1246
rect 708 1233 712 1242
rect 630 1228 648 1232
rect 655 1229 712 1233
rect 744 1232 748 1235
rect 552 1215 576 1219
rect 630 1215 634 1228
rect 655 1226 659 1229
rect 647 1218 651 1221
rect 558 1210 562 1215
rect 641 1214 665 1218
rect 558 1183 562 1186
rect 689 1185 693 1229
rect 738 1228 762 1232
rect 816 1229 820 1247
rect 833 1242 837 1247
rect 841 1231 845 1236
rect 854 1231 858 1253
rect 873 1240 877 1246
rect 816 1225 834 1229
rect 841 1227 858 1231
rect 738 1212 762 1216
rect 816 1212 820 1225
rect 841 1223 845 1227
rect 833 1215 837 1218
rect 744 1207 748 1212
rect 827 1211 851 1215
rect 854 1212 858 1227
rect 873 1218 877 1228
rect 942 1231 946 1250
rect 968 1231 972 1257
rect 942 1227 972 1231
rect 942 1223 946 1227
rect 873 1214 930 1218
rect 873 1213 877 1214
rect 854 1208 862 1212
rect 871 1197 891 1201
rect 552 1179 576 1183
rect 646 1181 693 1185
rect 470 1141 623 1145
rect 362 1123 420 1126
rect 263 1122 420 1123
rect 263 1119 366 1122
rect 491 1097 597 1100
rect 422 1096 597 1097
rect 422 1093 495 1096
rect 516 1095 597 1096
rect 516 1093 550 1095
rect 422 1092 426 1093
rect 389 1088 426 1092
rect 459 1091 495 1093
rect 405 1082 409 1088
rect 474 1086 478 1091
rect 531 1089 535 1093
rect 579 1089 583 1095
rect 500 1081 520 1085
rect 405 1064 409 1070
rect 405 1042 409 1052
rect 474 1055 478 1074
rect 500 1055 504 1081
rect 474 1051 504 1055
rect 474 1047 478 1051
rect 405 1038 462 1042
rect 405 1037 409 1038
rect 389 1021 423 1025
rect 419 1005 423 1021
rect 475 1022 479 1034
rect 500 1020 504 1051
rect 531 1058 535 1077
rect 587 1063 591 1083
rect 566 1059 580 1063
rect 587 1059 604 1063
rect 566 1058 570 1059
rect 531 1054 570 1058
rect 587 1056 591 1059
rect 531 1050 535 1054
rect 579 1041 583 1051
rect 532 1025 536 1037
rect 572 1037 583 1041
rect 500 1016 519 1020
rect 475 1005 479 1009
rect 532 1008 536 1012
rect 572 1008 576 1037
rect 518 1005 576 1008
rect 419 1004 576 1005
rect 419 1001 522 1004
rect 618 998 623 1141
rect 646 1091 650 1181
rect 657 1162 674 1166
rect 657 1134 661 1162
rect 681 1145 685 1169
rect 689 1166 693 1181
rect 744 1180 748 1183
rect 887 1181 891 1197
rect 943 1198 947 1210
rect 968 1196 972 1227
rect 999 1234 1003 1253
rect 1055 1239 1059 1259
rect 1232 1259 1236 1265
rect 1034 1235 1048 1239
rect 1055 1235 1065 1239
rect 1232 1237 1236 1247
rect 1273 1250 1277 1269
rect 1299 1250 1303 1276
rect 1273 1246 1303 1250
rect 1273 1242 1277 1246
rect 1034 1234 1038 1235
rect 999 1230 1038 1234
rect 1055 1232 1059 1235
rect 999 1226 1003 1230
rect 1232 1233 1261 1237
rect 1232 1232 1236 1233
rect 1047 1217 1051 1227
rect 1000 1201 1004 1213
rect 1040 1213 1051 1217
rect 1216 1216 1250 1220
rect 968 1192 987 1196
rect 943 1181 947 1185
rect 1000 1184 1004 1188
rect 1040 1184 1044 1213
rect 1246 1200 1250 1216
rect 1274 1217 1278 1229
rect 1299 1215 1303 1246
rect 1319 1253 1323 1272
rect 1359 1258 1363 1278
rect 1410 1269 1414 1296
rect 1419 1287 1443 1291
rect 1425 1282 1429 1287
rect 1480 1276 1484 1296
rect 1601 1293 1675 1298
rect 1808 1293 1887 1296
rect 1508 1270 1532 1274
rect 1384 1265 1426 1269
rect 1384 1258 1388 1265
rect 1338 1254 1352 1258
rect 1359 1254 1388 1258
rect 1338 1253 1342 1254
rect 1319 1249 1342 1253
rect 1359 1251 1363 1254
rect 1319 1245 1323 1249
rect 1351 1236 1355 1246
rect 1320 1220 1324 1232
rect 1344 1232 1355 1236
rect 1299 1211 1307 1215
rect 1274 1200 1278 1204
rect 1320 1203 1324 1207
rect 1344 1203 1348 1232
rect 1306 1200 1348 1203
rect 1246 1199 1348 1200
rect 1246 1196 1310 1199
rect 1313 1184 1392 1187
rect 986 1181 1044 1184
rect 887 1180 1044 1181
rect 1272 1183 1392 1184
rect 1272 1180 1317 1183
rect 1327 1182 1392 1183
rect 1327 1180 1361 1182
rect 738 1176 762 1180
rect 887 1177 990 1180
rect 1272 1179 1276 1180
rect 1239 1175 1276 1179
rect 1281 1178 1317 1180
rect 1255 1169 1259 1175
rect 1296 1173 1300 1178
rect 1342 1176 1346 1180
rect 1374 1176 1378 1182
rect 689 1162 700 1166
rect 1322 1168 1331 1172
rect 707 1145 711 1153
rect 1255 1151 1259 1157
rect 681 1141 711 1145
rect 662 1129 682 1133
rect 689 1126 693 1141
rect 1255 1129 1259 1139
rect 1296 1142 1300 1161
rect 1322 1142 1326 1168
rect 1296 1138 1326 1142
rect 1296 1134 1300 1138
rect 787 1124 834 1128
rect 681 1100 685 1120
rect 632 1087 682 1091
rect 647 1045 694 1049
rect 647 955 651 1045
rect 658 1026 675 1030
rect 658 998 662 1026
rect 682 1009 686 1033
rect 690 1030 694 1045
rect 787 1034 791 1124
rect 798 1105 815 1109
rect 798 1077 802 1105
rect 822 1088 826 1112
rect 830 1109 834 1124
rect 1255 1125 1284 1129
rect 1255 1124 1259 1125
rect 830 1105 841 1109
rect 1239 1108 1273 1112
rect 848 1088 852 1096
rect 1269 1092 1273 1108
rect 1297 1109 1301 1121
rect 1322 1107 1326 1138
rect 1342 1145 1346 1164
rect 1403 1163 1407 1265
rect 1425 1255 1429 1258
rect 1419 1251 1443 1255
rect 1497 1252 1501 1270
rect 1514 1265 1518 1270
rect 1601 1266 1605 1293
rect 1610 1284 1634 1288
rect 1616 1279 1620 1284
rect 1671 1273 1675 1293
rect 1767 1292 1887 1293
rect 1767 1289 1812 1292
rect 1822 1291 1887 1292
rect 1822 1289 1856 1291
rect 1767 1288 1771 1289
rect 1734 1284 1771 1288
rect 1776 1287 1812 1289
rect 1750 1278 1754 1284
rect 1791 1282 1795 1287
rect 1837 1285 1841 1289
rect 1869 1285 1873 1291
rect 1731 1273 1739 1277
rect 1817 1277 1826 1281
rect 1699 1267 1723 1271
rect 1522 1253 1526 1259
rect 1601 1262 1617 1266
rect 1601 1253 1605 1262
rect 1497 1248 1515 1252
rect 1522 1251 1605 1253
rect 1616 1252 1620 1255
rect 1522 1249 1551 1251
rect 1419 1235 1443 1239
rect 1497 1235 1501 1248
rect 1522 1246 1526 1249
rect 1556 1249 1605 1251
rect 1514 1238 1518 1241
rect 1425 1230 1429 1235
rect 1508 1234 1532 1238
rect 1425 1203 1429 1206
rect 1419 1199 1443 1203
rect 1592 1166 1597 1249
rect 1610 1248 1634 1252
rect 1688 1249 1692 1267
rect 1705 1262 1709 1267
rect 1713 1250 1717 1256
rect 1731 1250 1735 1273
rect 1750 1260 1754 1266
rect 1688 1245 1706 1249
rect 1713 1246 1735 1250
rect 1610 1232 1634 1236
rect 1688 1232 1692 1245
rect 1713 1243 1717 1246
rect 1705 1235 1709 1238
rect 1616 1227 1620 1232
rect 1699 1231 1723 1235
rect 1731 1232 1735 1246
rect 1750 1238 1754 1248
rect 1791 1251 1795 1270
rect 1817 1251 1821 1277
rect 1791 1247 1821 1251
rect 1791 1243 1795 1247
rect 1750 1234 1779 1238
rect 1750 1233 1754 1234
rect 1731 1228 1739 1232
rect 1734 1217 1768 1221
rect 1616 1200 1620 1203
rect 1764 1201 1768 1217
rect 1792 1218 1796 1230
rect 1817 1216 1821 1247
rect 1837 1254 1841 1273
rect 1877 1259 1881 1279
rect 1856 1255 1870 1259
rect 1877 1255 1887 1259
rect 1856 1254 1860 1255
rect 1837 1250 1860 1254
rect 1877 1252 1881 1255
rect 1837 1246 1841 1250
rect 1869 1237 1873 1247
rect 1838 1221 1842 1233
rect 1862 1233 1873 1237
rect 1817 1212 1825 1216
rect 1792 1201 1796 1205
rect 1838 1204 1842 1208
rect 1862 1204 1866 1233
rect 1824 1201 1866 1204
rect 1764 1200 1866 1201
rect 1610 1196 1634 1200
rect 1764 1197 1828 1200
rect 1403 1159 1450 1163
rect 1592 1162 1766 1166
rect 1361 1146 1375 1150
rect 1361 1145 1365 1146
rect 1342 1141 1365 1145
rect 1342 1137 1346 1141
rect 1374 1128 1378 1138
rect 1343 1112 1347 1124
rect 1367 1124 1378 1128
rect 1322 1103 1330 1107
rect 1297 1092 1301 1096
rect 1343 1095 1347 1099
rect 1367 1095 1371 1124
rect 1329 1092 1371 1095
rect 1269 1091 1371 1092
rect 1269 1088 1333 1091
rect 822 1084 852 1088
rect 803 1072 823 1076
rect 830 1069 834 1084
rect 1403 1069 1407 1159
rect 1414 1140 1431 1144
rect 1414 1112 1418 1140
rect 1438 1123 1442 1147
rect 1446 1144 1450 1159
rect 1539 1150 1579 1154
rect 1446 1140 1457 1144
rect 1539 1139 1543 1150
rect 1464 1123 1468 1131
rect 1438 1119 1468 1123
rect 1507 1135 1543 1139
rect 1419 1107 1439 1111
rect 1446 1104 1450 1119
rect 1438 1078 1442 1098
rect 1459 1092 1463 1119
rect 1469 1110 1493 1114
rect 1475 1105 1479 1110
rect 1483 1092 1487 1099
rect 1507 1092 1511 1135
rect 1459 1088 1476 1092
rect 1483 1088 1511 1092
rect 1483 1086 1487 1088
rect 1475 1078 1479 1081
rect 1469 1074 1493 1078
rect 1403 1065 1439 1069
rect 822 1043 826 1063
rect 1539 1050 1543 1135
rect 1578 1123 1582 1135
rect 1578 1119 1605 1123
rect 1578 1113 1582 1119
rect 1601 1113 1605 1119
rect 1570 1088 1574 1101
rect 1609 1088 1613 1101
rect 1625 1097 1649 1101
rect 1570 1084 1613 1088
rect 1631 1092 1635 1097
rect 1571 1059 1575 1084
rect 1602 1072 1606 1084
rect 1609 1079 1613 1084
rect 1609 1075 1632 1079
rect 1539 1046 1572 1050
rect 1594 1046 1598 1066
rect 1631 1065 1635 1068
rect 1625 1061 1649 1065
rect 1697 1049 1701 1162
rect 1708 1148 1746 1152
rect 1708 1058 1712 1148
rect 1718 1130 1727 1134
rect 1718 1097 1722 1130
rect 1734 1105 1738 1115
rect 1753 1105 1757 1133
rect 1773 1105 1777 1147
rect 1836 1151 1869 1155
rect 1799 1123 1823 1127
rect 1805 1118 1809 1123
rect 1813 1105 1817 1112
rect 1836 1105 1840 1151
rect 1848 1119 1869 1123
rect 1876 1116 1880 1136
rect 1895 1126 1919 1130
rect 1734 1101 1806 1105
rect 1813 1101 1840 1105
rect 1718 1093 1750 1097
rect 1757 1090 1761 1101
rect 1813 1099 1817 1101
rect 1805 1091 1809 1094
rect 1799 1087 1823 1091
rect 1749 1070 1753 1081
rect 1836 1070 1840 1101
rect 1901 1121 1905 1126
rect 1909 1109 1913 1115
rect 1886 1104 1902 1108
rect 1909 1105 1919 1109
rect 1868 1096 1872 1104
rect 1886 1096 1890 1104
rect 1909 1102 1913 1105
rect 1868 1092 1890 1096
rect 1901 1094 1905 1097
rect 1848 1082 1861 1086
rect 1868 1079 1872 1092
rect 1878 1086 1882 1092
rect 1895 1090 1919 1094
rect 1879 1070 1883 1073
rect 1836 1066 1883 1070
rect 1708 1054 1750 1058
rect 1697 1045 1750 1049
rect 1757 1042 1761 1061
rect 787 1030 823 1034
rect 690 1026 701 1030
rect 708 1009 712 1017
rect 787 1009 790 1030
rect 682 1005 790 1009
rect 663 993 683 997
rect 690 990 694 1005
rect 682 964 686 984
rect 633 951 683 955
rect 818 913 924 916
rect 772 912 924 913
rect 772 909 822 912
rect 843 911 924 912
rect 843 909 877 911
rect 772 908 776 909
rect 739 904 776 908
rect 786 907 822 909
rect 755 898 759 904
rect 801 902 805 907
rect 858 905 862 909
rect 906 905 910 911
rect 944 906 1018 911
rect 827 897 847 901
rect 755 880 759 886
rect 755 858 759 868
rect 801 871 805 890
rect 827 871 831 897
rect 801 867 831 871
rect 801 863 805 867
rect 755 854 789 858
rect 755 853 759 854
rect 739 837 773 841
rect 769 821 773 837
rect 802 838 806 850
rect 827 836 831 867
rect 858 874 862 893
rect 914 879 918 899
rect 944 879 948 906
rect 953 897 977 901
rect 959 892 963 897
rect 1014 886 1018 906
rect 1105 903 1179 908
rect 1042 880 1066 884
rect 893 875 907 879
rect 914 875 960 879
rect 893 874 897 875
rect 858 870 897 874
rect 914 872 918 875
rect 858 866 862 870
rect 906 857 910 867
rect 859 841 863 853
rect 899 853 910 857
rect 827 832 846 836
rect 802 821 806 825
rect 859 824 863 828
rect 899 824 903 853
rect 845 821 903 824
rect 769 820 903 821
rect 769 817 849 820
rect 843 782 928 785
rect 802 781 928 782
rect 802 778 847 781
rect 860 780 928 781
rect 860 778 894 780
rect 802 777 806 778
rect 769 773 806 777
rect 811 776 847 778
rect 785 767 789 773
rect 826 771 830 776
rect 875 774 879 778
rect 910 774 914 780
rect 937 775 941 875
rect 959 865 963 868
rect 953 861 977 865
rect 1031 862 1035 880
rect 1048 875 1052 880
rect 1105 876 1109 903
rect 1114 894 1138 898
rect 1120 889 1124 894
rect 1175 883 1179 903
rect 1326 889 1422 892
rect 1281 888 1422 889
rect 1281 885 1330 888
rect 1351 887 1422 888
rect 1351 885 1385 887
rect 1281 884 1285 885
rect 1203 877 1227 881
rect 1248 880 1285 884
rect 1294 883 1330 885
rect 1056 863 1060 869
rect 1084 872 1121 876
rect 1084 865 1090 872
rect 1031 858 1049 862
rect 1056 859 1084 863
rect 1120 862 1124 865
rect 953 845 977 849
rect 1031 845 1035 858
rect 1056 856 1060 859
rect 1114 858 1138 862
rect 1192 859 1196 877
rect 1209 872 1213 877
rect 1264 874 1268 880
rect 1309 878 1313 883
rect 1366 881 1370 885
rect 1404 881 1408 887
rect 1217 860 1221 866
rect 1233 869 1253 873
rect 1335 873 1355 877
rect 1233 860 1237 869
rect 1192 855 1210 859
rect 1217 856 1237 860
rect 1048 848 1052 851
rect 959 840 963 845
rect 1042 844 1066 848
rect 1114 842 1138 846
rect 1192 842 1196 855
rect 1217 853 1221 856
rect 1209 845 1213 848
rect 1120 837 1124 842
rect 1203 841 1227 845
rect 1233 828 1237 856
rect 1264 856 1268 862
rect 1264 834 1268 844
rect 1309 847 1313 866
rect 1335 847 1339 873
rect 1309 843 1339 847
rect 1309 839 1313 843
rect 1264 830 1297 834
rect 1264 829 1268 830
rect 1233 824 1253 828
rect 959 813 963 816
rect 1248 813 1282 817
rect 953 809 977 813
rect 1120 810 1124 813
rect 1114 806 1138 810
rect 1278 797 1282 813
rect 1310 814 1314 826
rect 1335 812 1339 843
rect 1366 850 1370 869
rect 1412 855 1416 875
rect 1391 851 1405 855
rect 1412 851 1422 855
rect 1391 850 1395 851
rect 1366 846 1395 850
rect 1412 848 1416 851
rect 1366 842 1370 846
rect 1735 843 1814 846
rect 1404 833 1408 843
rect 1694 842 1814 843
rect 1694 839 1739 842
rect 1749 841 1814 842
rect 1749 839 1783 841
rect 1694 838 1698 839
rect 1661 834 1698 838
rect 1703 837 1739 839
rect 1367 817 1371 829
rect 1397 829 1408 833
rect 1335 808 1354 812
rect 1310 797 1314 801
rect 1367 800 1371 804
rect 1397 800 1401 829
rect 1677 828 1681 834
rect 1718 832 1722 837
rect 1764 835 1768 839
rect 1796 835 1800 841
rect 1832 836 1906 841
rect 1744 827 1753 831
rect 1677 810 1681 816
rect 1353 797 1401 800
rect 1278 796 1401 797
rect 1278 793 1357 796
rect 1677 788 1681 798
rect 1718 801 1722 820
rect 1744 801 1748 827
rect 1718 797 1748 801
rect 1718 793 1722 797
rect 1677 784 1706 788
rect 1677 783 1681 784
rect 852 766 864 770
rect 937 771 984 775
rect 785 749 789 755
rect 785 727 789 737
rect 826 740 830 759
rect 852 740 856 766
rect 826 736 856 740
rect 826 732 830 736
rect 785 723 814 727
rect 785 722 789 723
rect 769 706 803 710
rect 799 690 803 706
rect 827 707 831 719
rect 852 705 856 736
rect 875 743 879 762
rect 897 744 911 748
rect 897 743 901 744
rect 875 739 901 743
rect 875 735 879 739
rect 910 726 914 736
rect 876 710 880 722
rect 903 722 914 726
rect 852 701 863 705
rect 827 690 831 694
rect 876 693 880 697
rect 903 693 907 722
rect 862 690 907 693
rect 799 689 907 690
rect 799 686 866 689
rect 937 681 941 771
rect 948 752 965 756
rect 948 724 952 752
rect 972 735 976 759
rect 980 756 984 771
rect 1073 774 1113 778
rect 980 752 991 756
rect 998 735 1002 743
rect 972 731 1002 735
rect 953 719 973 723
rect 980 716 984 731
rect 972 690 976 710
rect 993 704 997 731
rect 1003 722 1027 726
rect 1009 717 1013 722
rect 1017 704 1021 711
rect 1073 704 1077 774
rect 1661 767 1695 771
rect 1112 747 1116 759
rect 1691 751 1695 767
rect 1719 768 1723 780
rect 1744 766 1748 797
rect 1764 804 1768 823
rect 1804 809 1808 829
rect 1832 809 1836 836
rect 1841 827 1865 831
rect 1847 822 1851 827
rect 1902 816 1906 836
rect 2092 833 2166 838
rect 1930 810 1954 814
rect 1783 805 1797 809
rect 1804 805 1848 809
rect 1783 804 1787 805
rect 1764 800 1787 804
rect 1804 802 1808 805
rect 1764 796 1768 800
rect 1796 787 1800 797
rect 1765 771 1769 783
rect 1789 783 1800 787
rect 1744 762 1752 766
rect 1719 751 1723 755
rect 1765 754 1769 758
rect 1789 754 1793 783
rect 1751 751 1793 754
rect 1691 750 1793 751
rect 1691 747 1755 750
rect 1112 743 1139 747
rect 1112 737 1116 743
rect 1135 737 1139 743
rect 1104 712 1108 725
rect 1143 712 1147 725
rect 1159 721 1183 725
rect 1104 708 1147 712
rect 1165 716 1169 721
rect 993 700 1010 704
rect 1017 700 1077 704
rect 1017 698 1021 700
rect 1009 690 1013 693
rect 1003 686 1027 690
rect 937 677 973 681
rect 1073 674 1077 700
rect 1105 683 1109 708
rect 1136 696 1140 708
rect 1143 703 1147 708
rect 1143 699 1166 703
rect 1735 701 1814 704
rect 1694 700 1814 701
rect 1694 697 1739 700
rect 1749 699 1814 700
rect 1749 697 1783 699
rect 1694 696 1698 697
rect 1661 692 1698 696
rect 1703 695 1739 697
rect 1073 670 1106 674
rect 1128 670 1132 690
rect 1165 689 1169 692
rect 1159 685 1183 689
rect 1677 686 1681 692
rect 1718 690 1722 695
rect 1764 693 1768 697
rect 1796 693 1800 699
rect 1744 685 1753 689
rect 1677 668 1681 674
rect 1677 646 1681 656
rect 1718 659 1722 678
rect 1744 659 1748 685
rect 1718 655 1748 659
rect 1718 651 1722 655
rect 1677 642 1706 646
rect 1677 641 1681 642
rect 1661 625 1695 629
rect 1691 609 1695 625
rect 1719 626 1723 638
rect 1744 624 1748 655
rect 1764 662 1768 681
rect 1783 663 1797 667
rect 1783 662 1787 663
rect 1764 658 1787 662
rect 1764 654 1768 658
rect 1796 645 1800 655
rect 1765 629 1769 641
rect 1789 641 1800 645
rect 1825 644 1829 805
rect 1847 795 1851 798
rect 1841 791 1865 795
rect 1919 792 1923 810
rect 1936 805 1940 810
rect 2092 806 2096 833
rect 2101 824 2125 828
rect 2107 819 2111 824
rect 2162 813 2166 833
rect 2299 823 2378 826
rect 2258 822 2378 823
rect 2258 819 2303 822
rect 2313 821 2378 822
rect 2313 819 2347 821
rect 2258 818 2262 819
rect 2225 814 2262 818
rect 2267 817 2303 819
rect 2190 807 2214 811
rect 2241 808 2245 814
rect 2282 812 2286 817
rect 2328 815 2332 819
rect 2360 815 2364 821
rect 1944 793 1948 799
rect 2071 802 2108 806
rect 2071 793 2075 802
rect 1919 788 1937 792
rect 1944 789 2075 793
rect 2107 792 2111 795
rect 1841 775 1865 779
rect 1919 775 1923 788
rect 1944 786 1948 789
rect 1936 778 1940 781
rect 1847 770 1851 775
rect 1930 774 1954 778
rect 1847 743 1851 746
rect 1841 739 1865 743
rect 1989 700 1993 789
rect 2065 724 2069 789
rect 2101 788 2125 792
rect 2179 789 2183 807
rect 2196 802 2200 807
rect 2220 803 2230 807
rect 2308 807 2317 811
rect 2204 790 2208 796
rect 2220 790 2224 803
rect 2179 785 2197 789
rect 2204 786 2224 790
rect 2241 790 2245 796
rect 2101 772 2125 776
rect 2179 772 2183 785
rect 2204 783 2208 786
rect 2196 775 2200 778
rect 2107 767 2111 772
rect 2190 771 2214 775
rect 2220 762 2224 786
rect 2241 768 2245 778
rect 2282 781 2286 800
rect 2308 781 2312 807
rect 2282 777 2312 781
rect 2282 773 2286 777
rect 2241 764 2270 768
rect 2241 763 2245 764
rect 2220 758 2230 762
rect 2225 747 2259 751
rect 2107 740 2111 743
rect 2101 736 2125 740
rect 2255 731 2259 747
rect 2283 748 2287 760
rect 2308 746 2312 777
rect 2328 784 2332 803
rect 2368 789 2372 809
rect 2347 785 2361 789
rect 2368 785 2378 789
rect 2347 784 2351 785
rect 2328 780 2351 784
rect 2368 782 2372 785
rect 2328 776 2332 780
rect 2360 767 2364 777
rect 2329 751 2333 763
rect 2353 763 2364 767
rect 2308 742 2316 746
rect 2283 731 2287 735
rect 2329 734 2333 738
rect 2353 734 2357 763
rect 2315 731 2357 734
rect 2255 730 2357 731
rect 2255 727 2319 730
rect 2065 719 2165 724
rect 1989 696 2087 700
rect 1744 620 1752 624
rect 1719 609 1723 613
rect 1765 612 1769 616
rect 1789 612 1793 641
rect 1751 609 1793 612
rect 1691 608 1793 609
rect 1825 640 1872 644
rect 1691 605 1755 608
rect 1825 550 1829 640
rect 1836 621 1853 625
rect 1836 593 1840 621
rect 1860 604 1864 628
rect 1868 625 1872 640
rect 1868 621 1879 625
rect 1886 604 1890 612
rect 1860 600 1890 604
rect 1841 588 1861 592
rect 1868 585 1872 600
rect 1860 559 1864 579
rect 1881 573 1885 600
rect 1895 591 1919 595
rect 1901 586 1905 591
rect 1909 573 1913 580
rect 1881 569 1902 573
rect 1909 569 1921 573
rect 1909 567 1913 569
rect 1901 559 1905 562
rect 1895 555 1919 559
rect 1825 546 1861 550
rect 1989 524 1993 696
rect 2265 684 2346 688
rect 2001 676 2070 680
rect 2001 563 2005 676
rect 2012 662 2050 666
rect 2012 572 2016 662
rect 2022 644 2031 648
rect 2022 611 2026 644
rect 2038 619 2042 629
rect 2057 619 2061 647
rect 2077 619 2081 661
rect 2094 619 2098 681
rect 2038 615 2098 619
rect 2148 672 2188 676
rect 2022 607 2054 611
rect 2061 604 2065 615
rect 2053 584 2057 595
rect 2012 568 2054 572
rect 2001 559 2054 563
rect 2061 556 2065 575
rect 2053 536 2057 547
rect 1989 520 2054 524
rect 2087 516 2094 615
rect 2148 602 2152 672
rect 2187 645 2191 657
rect 2187 641 2214 645
rect 2187 635 2191 641
rect 2210 635 2214 641
rect 2179 610 2183 623
rect 2218 610 2222 623
rect 2234 619 2258 623
rect 2179 606 2222 610
rect 2240 614 2244 619
rect 2136 598 2152 602
rect 2148 572 2152 598
rect 2180 581 2184 606
rect 2211 594 2215 606
rect 2218 601 2222 606
rect 2218 597 2241 601
rect 2148 568 2181 572
rect 2203 568 2207 588
rect 2240 587 2244 590
rect 2234 583 2258 587
rect 2277 571 2281 684
rect 2288 670 2326 674
rect 2288 580 2292 670
rect 2714 679 2793 682
rect 2673 678 2793 679
rect 2298 652 2307 656
rect 2298 619 2302 652
rect 2314 627 2318 637
rect 2333 627 2337 655
rect 2353 627 2357 669
rect 2408 673 2441 677
rect 2522 673 2570 677
rect 2673 675 2718 678
rect 2728 677 2793 678
rect 2728 675 2762 677
rect 2673 674 2677 675
rect 2375 645 2399 649
rect 2381 640 2385 645
rect 2389 627 2393 634
rect 2408 627 2412 673
rect 2420 641 2441 645
rect 2448 638 2452 658
rect 2314 623 2382 627
rect 2389 623 2412 627
rect 2298 615 2330 619
rect 2337 612 2341 623
rect 2389 621 2393 623
rect 2381 613 2385 616
rect 2375 609 2399 613
rect 2329 592 2333 603
rect 2408 592 2412 623
rect 2479 636 2503 640
rect 2485 631 2489 636
rect 2440 618 2444 626
rect 2493 618 2497 625
rect 2522 618 2526 673
rect 2640 670 2677 674
rect 2682 673 2718 675
rect 2656 664 2660 670
rect 2697 668 2701 673
rect 2743 671 2747 675
rect 2775 671 2779 677
rect 2539 641 2570 645
rect 2440 614 2486 618
rect 2493 614 2529 618
rect 2420 604 2433 608
rect 2440 601 2444 614
rect 2450 608 2454 614
rect 2493 612 2497 614
rect 2525 609 2529 614
rect 2485 604 2489 607
rect 2479 600 2503 604
rect 2451 592 2455 595
rect 2408 588 2455 592
rect 2539 592 2543 641
rect 2577 638 2581 658
rect 2630 659 2645 663
rect 2723 663 2732 667
rect 2597 636 2621 640
rect 2603 631 2607 636
rect 2569 618 2573 626
rect 2611 618 2615 625
rect 2630 618 2634 659
rect 2656 646 2660 652
rect 2656 624 2660 634
rect 2697 637 2701 656
rect 2723 637 2727 663
rect 2697 633 2727 637
rect 2697 629 2701 633
rect 2656 620 2685 624
rect 2656 619 2660 620
rect 2569 614 2604 618
rect 2611 614 2645 618
rect 2569 601 2573 614
rect 2579 608 2583 614
rect 2611 612 2615 614
rect 2603 604 2607 607
rect 2597 600 2621 604
rect 2640 603 2674 607
rect 2580 592 2584 595
rect 2539 588 2584 592
rect 2288 576 2330 580
rect 2277 567 2330 571
rect 2337 564 2341 583
rect 2107 533 2131 537
rect 2113 528 2117 533
rect 2087 515 2103 516
rect 2121 515 2125 522
rect 2539 516 2544 588
rect 2670 587 2674 603
rect 2698 604 2702 616
rect 2723 602 2727 633
rect 2743 640 2747 659
rect 2783 645 2787 665
rect 2762 641 2776 645
rect 2783 641 2793 645
rect 2762 640 2766 641
rect 2743 636 2766 640
rect 2783 638 2787 641
rect 2743 632 2747 636
rect 2775 623 2779 633
rect 2744 607 2748 619
rect 2768 619 2779 623
rect 2723 598 2731 602
rect 2698 587 2702 591
rect 2744 590 2748 594
rect 2768 590 2772 619
rect 2730 587 2772 590
rect 2670 586 2772 587
rect 2670 583 2734 586
rect 2134 515 2544 516
rect 2087 511 2114 515
rect 2121 511 2544 515
rect 2087 510 2103 511
rect 2121 509 2125 511
rect 2134 510 2544 511
rect 2113 501 2117 504
rect 2107 497 2131 501
<< m2contact >>
rect 438 1177 443 1182
rect 604 1059 609 1064
rect 657 1129 662 1134
rect 706 1136 711 1141
rect 618 993 623 998
rect 798 1072 803 1077
rect 1414 1107 1419 1112
rect 658 993 663 998
rect 948 719 953 724
rect 1836 588 1841 593
rect 2525 604 2530 609
<< metal2 >>
rect 1473 1261 1485 1266
rect 1473 1246 1477 1261
rect 1664 1258 1676 1263
rect 606 1241 618 1246
rect 606 1226 610 1241
rect 544 1222 610 1226
rect 792 1238 804 1243
rect 1411 1242 1477 1246
rect 1664 1243 1668 1258
rect 792 1223 796 1238
rect 544 1200 548 1222
rect 730 1219 796 1223
rect 1411 1220 1415 1242
rect 1602 1239 1668 1243
rect 517 1197 548 1200
rect 566 1197 570 1204
rect 609 1200 618 1204
rect 609 1197 613 1200
rect 730 1197 734 1219
rect 1396 1217 1415 1220
rect 1433 1217 1437 1224
rect 1476 1220 1485 1224
rect 1476 1217 1480 1220
rect 1396 1216 1425 1217
rect 517 1196 558 1197
rect 517 1181 521 1196
rect 544 1193 558 1196
rect 566 1193 613 1197
rect 640 1194 734 1197
rect 752 1194 756 1201
rect 795 1197 804 1201
rect 795 1194 799 1197
rect 640 1193 744 1194
rect 566 1191 570 1193
rect 443 1177 521 1181
rect 640 1134 644 1193
rect 730 1190 744 1193
rect 752 1190 799 1194
rect 752 1188 756 1190
rect 1382 1154 1386 1170
rect 1396 1154 1400 1216
rect 1411 1213 1425 1216
rect 1433 1213 1480 1217
rect 1602 1214 1606 1239
rect 1624 1214 1628 1221
rect 1667 1217 1676 1221
rect 1667 1214 1671 1217
rect 1433 1211 1437 1213
rect 1602 1210 1616 1214
rect 1624 1210 1671 1214
rect 1624 1208 1628 1210
rect 1382 1150 1400 1154
rect 1382 1143 1386 1150
rect 604 1129 657 1134
rect 604 1064 609 1129
rect 707 1077 711 1136
rect 1396 1112 1400 1150
rect 1396 1107 1414 1112
rect 1591 1094 1602 1098
rect 1591 1084 1595 1094
rect 1563 1080 1595 1084
rect 707 1072 798 1077
rect 1591 1075 1595 1080
rect 623 993 658 998
rect 1007 871 1019 876
rect 1007 856 1011 871
rect 1168 868 1180 873
rect 945 852 1011 856
rect 1168 853 1172 868
rect 945 830 949 852
rect 1106 849 1172 853
rect 930 827 949 830
rect 967 827 971 834
rect 1010 830 1019 834
rect 1010 827 1014 830
rect 1106 827 1110 849
rect 930 826 959 827
rect 918 750 922 768
rect 930 750 934 826
rect 945 823 959 826
rect 967 823 1014 827
rect 1083 824 1110 827
rect 1128 824 1132 831
rect 1171 827 1180 831
rect 1171 824 1175 827
rect 1083 823 1120 824
rect 967 821 971 823
rect 918 746 934 750
rect 918 741 922 746
rect 930 724 934 746
rect 930 719 948 724
rect 1083 708 1087 823
rect 1106 820 1120 823
rect 1128 820 1175 824
rect 1128 818 1132 820
rect 1895 801 1907 806
rect 1895 786 1899 801
rect 1833 782 1899 786
rect 2155 798 2167 803
rect 2155 783 2159 798
rect 1833 760 1837 782
rect 2093 779 2159 783
rect 1818 757 1837 760
rect 1855 757 1859 764
rect 1898 760 1907 764
rect 1898 757 1902 760
rect 2093 757 2097 779
rect 1818 756 1847 757
rect 1125 718 1136 722
rect 1125 708 1129 718
rect 1083 704 1129 708
rect 1125 699 1129 704
rect 1804 669 1808 687
rect 1818 669 1822 756
rect 1833 753 1847 756
rect 1855 753 1902 757
rect 1980 754 2097 757
rect 2115 754 2119 761
rect 2158 757 2167 761
rect 2158 754 2162 757
rect 1980 753 2107 754
rect 1855 751 1859 753
rect 2093 750 2107 753
rect 2115 750 2162 754
rect 2115 748 2119 750
rect 1804 665 1822 669
rect 1804 660 1808 665
rect 1818 593 1822 665
rect 2200 616 2211 620
rect 2200 606 2204 616
rect 2172 602 2204 606
rect 2530 604 2562 608
rect 2200 597 2204 602
rect 1818 588 1836 593
<< m3contact >>
rect 2160 719 2165 724
<< m123contact >>
rect 1551 1245 1556 1251
rect 1843 1118 1848 1123
rect 1843 1081 1848 1086
rect 1084 859 1090 865
rect 2415 640 2420 645
rect 2415 603 2420 608
<< metal3 >>
rect 1433 1270 1437 1276
rect 1433 1265 1465 1270
rect 1433 1263 1437 1265
rect 566 1250 570 1256
rect 566 1245 598 1250
rect 566 1243 570 1245
rect 594 1215 598 1245
rect 752 1247 756 1253
rect 752 1242 784 1247
rect 752 1240 756 1242
rect 594 1209 613 1215
rect 780 1212 784 1242
rect 1461 1235 1465 1265
rect 1624 1267 1628 1273
rect 1624 1262 1656 1267
rect 1624 1260 1628 1262
rect 1461 1229 1480 1235
rect 780 1206 799 1212
rect 1551 1120 1555 1245
rect 1652 1232 1656 1262
rect 1652 1226 1671 1232
rect 1551 1116 1571 1120
rect 1551 1037 1555 1116
rect 1843 1086 1848 1118
rect 1639 1079 1643 1086
rect 1639 1075 1670 1079
rect 1639 1073 1643 1075
rect 1551 1033 1595 1037
rect 1666 1027 1670 1075
rect 1843 1027 1848 1081
rect 1666 1023 1848 1027
rect 967 880 971 886
rect 967 875 999 880
rect 967 873 971 875
rect 995 845 999 875
rect 1128 877 1132 883
rect 1128 872 1160 877
rect 1128 870 1132 872
rect 995 839 1014 845
rect 1085 744 1089 859
rect 1156 842 1160 872
rect 1156 836 1175 842
rect 1855 810 1859 816
rect 1855 805 1887 810
rect 1855 803 1859 805
rect 1883 775 1887 805
rect 2115 807 2119 813
rect 2115 802 2147 807
rect 2115 800 2119 802
rect 1883 769 1902 775
rect 2143 772 2147 802
rect 2143 766 2162 772
rect 1085 740 1105 744
rect 1085 661 1089 740
rect 1173 703 1177 710
rect 1173 699 1183 703
rect 1173 697 1177 699
rect 1085 657 1129 661
rect 2160 642 2164 719
rect 2160 638 2180 642
rect 2160 559 2164 638
rect 2415 608 2420 640
rect 2248 601 2252 608
rect 2248 597 2279 601
rect 2248 595 2252 597
rect 2160 555 2204 559
rect 2275 549 2279 597
rect 2415 549 2420 603
rect 2275 545 2420 549
<< labels >>
rlabel nwell 572 1264 574 1266 1 vdd
rlabel pdcontact 558 1256 562 1262 1 vdd
rlabel nwell 572 1212 574 1214 1 vdd
rlabel pdcontact 558 1204 562 1210 1 vdd
rlabel nwell 661 1247 663 1249 1 vdd
rlabel pdcontact 647 1239 651 1245 1 vdd
rlabel ndcontact 647 1221 651 1225 1 gnd
rlabel ndcontact 558 1238 562 1242 1 gnd
rlabel ndcontact 558 1186 562 1190 1 gnd
rlabel polycontact 559 1245 563 1249 1 A0
rlabel ndcontact 566 1239 570 1243 1 A0N1
rlabel pdcontact 566 1256 570 1262 1 A0N1
rlabel polycontact 558 1193 562 1197 1 B0
rlabel ndcontact 566 1187 570 1191 1 B0N1
rlabel pdcontact 566 1204 570 1210 1 B0N1
rlabel polycontact 618 1200 622 1204 1 B0N1
rlabel ndcontact 613 1209 617 1214 1 A0N1
rlabel polycontact 618 1241 622 1246 1 B0
rlabel ndcontact 613 1250 617 1255 1 A0
rlabel ndcontact 630 1251 634 1255 1 X0
rlabel ndcontact 630 1210 634 1214 1 X0
rlabel polycontact 648 1228 652 1232 1 X0
rlabel pdcontact 655 1239 659 1245 1 P0
rlabel ndcontact 655 1222 659 1226 1 P0
rlabel pdcontact 699 1153 703 1159 1 vdd
rlabel pdcontact 673 1169 677 1175 1 vdd
rlabel ndcontact 689 1094 693 1100 1 gnd
rlabel pdcontact 700 1017 704 1023 1 vdd
rlabel pdcontact 674 1033 678 1039 1 vdd
rlabel ndcontact 690 958 694 964 1 gnd
rlabel pdcontact 840 1096 844 1102 1 vdd
rlabel pdcontact 814 1112 818 1118 1 vdd
rlabel ndcontact 830 1037 834 1043 1 gnd
rlabel m2contact 658 993 662 997 1 A0
rlabel polycontact 683 993 687 997 1 A0
rlabel polycontact 675 1026 679 1030 1 A0
rlabel polycontact 683 951 687 955 1 B0
rlabel polycontact 701 1026 705 1030 1 B0
rlabel pdcontact 682 1034 686 1038 1 Y0
rlabel pdcontact 708 1018 712 1022 1 Y0
rlabel ndcontact 690 985 694 989 1 Y0
rlabel ndcontact 682 985 686 989 1 N0
rlabel ndcontact 682 959 686 963 1 N0
rlabel polycontact 682 1087 686 1091 1 P0
rlabel polycontact 700 1162 704 1166 1 P0
rlabel m2contact 657 1129 661 1133 1 C0
rlabel polycontact 682 1129 686 1133 1 C0
rlabel polycontact 674 1162 678 1166 1 C0
rlabel pdcontact 681 1170 685 1174 1 Z0
rlabel pdcontact 707 1154 711 1158 1 Z0
rlabel ndcontact 689 1121 693 1125 1 Z0
rlabel ndcontact 681 1121 685 1125 1 M0
rlabel ndcontact 681 1095 685 1099 1 M0
rlabel m2contact 708 1137 710 1139 1 Z0
rlabel m2contact 798 1072 802 1076 1 Z0
rlabel polycontact 823 1072 827 1076 1 Z0
rlabel polycontact 815 1105 819 1109 1 Z0
rlabel polycontact 823 1030 827 1034 1 Y0
rlabel polycontact 841 1105 845 1109 1 Y0
rlabel ndcontact 822 1064 826 1068 1 K0
rlabel ndcontact 822 1038 826 1042 1 K0
rlabel pdcontact 848 1096 852 1100 1 C1
rlabel pdcontact 822 1113 826 1117 1 C1
rlabel ndcontact 830 1064 834 1068 1 C1
rlabel nwell 698 1174 702 1178 1 vdd
rlabel nwell 842 1115 846 1119 1 vdd
rlabel nwell 707 1035 711 1039 1 vdd
rlabel polycontact 245 1286 249 1290 1 clk
rlabel polycontact 313 1240 317 1244 1 clk
rlabel polycontact 314 1305 318 1309 1 clk
rlabel polycontact 370 1268 374 1272 1 clk
rlabel metal1 314 1320 339 1324 1 vdd
rlabel metal1 373 1323 398 1327 5 vdd
rlabel metal1 422 1322 447 1326 5 vdd
rlabel metal1 367 1320 401 1324 1 vdd
rlabel metal1 310 1318 344 1322 1 vdd
rlabel metal1 240 1315 276 1319 5 vdd
rlabel metal1 240 1315 276 1318 1 vdd
rlabel metal1 423 1322 448 1324 5 vdd
rlabel nwell 389 1314 392 1317 1 vdd
rlabel nwell 332 1311 335 1314 1 vdd
rlabel nwell 270 1310 273 1313 1 vdd
rlabel nwell 444 1317 447 1320 7 vdd
rlabel pdcontact 256 1305 260 1309 1 vdd
rlabel ndcontact 256 1252 260 1256 1 gnd
rlabel ndcontact 326 1236 330 1240 1 gnd
rlabel ndcontact 383 1239 387 1243 1 gnd
rlabel ndcontact 430 1278 434 1282 1 gnd
rlabel pdcontact 325 1309 329 1313 1 vdd
rlabel pdcontact 382 1312 386 1316 1 vdd
rlabel pdcontact 430 1310 434 1316 1 vdd
rlabel ndcontact 438 1279 442 1283 1 A0
rlabel pdcontact 438 1310 442 1314 1 A0
rlabel polycontact 245 1259 249 1263 1 AA0
rlabel polycontact 245 1304 249 1308 1 AA0
rlabel pdcontact 256 1297 260 1301 1 AV1
rlabel pdcontact 256 1287 260 1291 1 AV1
rlabel pdcontact 256 1279 260 1283 1 AV2
rlabel ndcontact 256 1260 260 1264 1 AV2
rlabel polycontact 313 1265 317 1269 1 AV2
rlabel ndcontact 326 1245 330 1249 1 AV3
rlabel ndcontact 326 1261 330 1265 1 AV3
rlabel ndcontact 325 1270 329 1274 1 AV4
rlabel pdcontact 325 1301 329 1305 1 AV4
rlabel polycontact 371 1308 375 1312 1 AV4
rlabel polycontact 370 1243 374 1247 1 AV4
rlabel ndcontact 383 1248 387 1252 1 AV5
rlabel ndcontact 383 1264 387 1268 1 AV5
rlabel ndcontact 382 1273 386 1277 1 AV6
rlabel pdcontact 382 1304 386 1308 1 AV6
rlabel polycontact 431 1286 435 1290 1 AV6
rlabel polycontact 238 1177 242 1181 1 clk
rlabel polycontact 306 1131 310 1135 1 clk
rlabel polycontact 307 1196 311 1200 1 clk
rlabel polycontact 363 1159 367 1163 1 clk
rlabel metal1 307 1211 332 1215 1 vdd
rlabel metal1 366 1214 391 1218 5 vdd
rlabel metal1 415 1213 440 1217 5 vdd
rlabel metal1 360 1211 394 1215 1 vdd
rlabel metal1 303 1209 337 1213 1 vdd
rlabel metal1 233 1206 269 1210 5 vdd
rlabel metal1 233 1206 269 1209 1 vdd
rlabel metal1 416 1213 441 1215 5 vdd
rlabel nwell 382 1205 385 1208 1 vdd
rlabel nwell 325 1202 328 1205 1 vdd
rlabel nwell 263 1201 266 1204 1 vdd
rlabel nwell 437 1208 440 1211 7 vdd
rlabel pdcontact 249 1196 253 1200 1 vdd
rlabel ndcontact 249 1143 253 1147 1 gnd
rlabel ndcontact 319 1127 323 1131 1 gnd
rlabel ndcontact 376 1130 380 1134 1 gnd
rlabel ndcontact 423 1169 427 1173 1 gnd
rlabel pdcontact 318 1200 322 1204 1 vdd
rlabel pdcontact 375 1203 379 1207 1 vdd
rlabel pdcontact 423 1201 427 1207 1 vdd
rlabel m2contact 439 1178 441 1180 1 B0
rlabel ndcontact 431 1170 435 1174 1 B0
rlabel pdcontact 431 1202 435 1206 1 B0
rlabel polycontact 238 1195 242 1199 1 BB0
rlabel polycontact 238 1150 242 1154 1 BB0
rlabel ndcontact 249 1151 253 1155 1 BY0
rlabel pdcontact 249 1170 253 1174 1 BY0
rlabel polycontact 306 1156 310 1160 1 BY0
rlabel pdcontact 249 1178 253 1182 1 BY1
rlabel pdcontact 249 1188 253 1192 1 BY1
rlabel ndcontact 319 1136 323 1140 1 BY2
rlabel ndcontact 319 1152 323 1156 1 BY2
rlabel ndcontact 318 1161 322 1165 1 BY3
rlabel pdcontact 318 1192 322 1196 1 BY3
rlabel polycontact 364 1199 368 1203 1 BY3
rlabel polycontact 363 1134 367 1138 1 BY3
rlabel ndcontact 376 1139 380 1143 1 BY4
rlabel ndcontact 376 1155 380 1159 1 BY4
rlabel ndcontact 375 1164 379 1168 1 BY5
rlabel pdcontact 375 1195 379 1199 1 BY5
rlabel polycontact 424 1177 428 1181 1 BY5
rlabel polycontact 394 1059 398 1063 1 clk
rlabel polycontact 462 1013 466 1017 1 clk
rlabel polycontact 463 1078 467 1082 1 clk
rlabel polycontact 519 1041 523 1045 1 clk
rlabel metal1 463 1093 488 1097 1 vdd
rlabel metal1 522 1096 547 1100 5 vdd
rlabel metal1 571 1095 596 1099 5 vdd
rlabel metal1 516 1093 550 1097 1 vdd
rlabel metal1 459 1091 493 1095 1 vdd
rlabel metal1 389 1088 425 1092 5 vdd
rlabel metal1 389 1088 425 1091 1 vdd
rlabel metal1 572 1095 597 1097 5 vdd
rlabel nwell 538 1087 541 1090 1 vdd
rlabel nwell 481 1084 484 1087 1 vdd
rlabel nwell 419 1083 422 1086 1 vdd
rlabel nwell 593 1090 596 1093 7 vdd
rlabel pdcontact 405 1078 409 1082 1 vdd
rlabel ndcontact 405 1025 409 1029 1 gnd
rlabel ndcontact 475 1009 479 1013 1 gnd
rlabel ndcontact 532 1012 536 1016 1 gnd
rlabel ndcontact 579 1051 583 1055 1 gnd
rlabel pdcontact 474 1082 478 1086 1 vdd
rlabel pdcontact 531 1085 535 1089 1 vdd
rlabel pdcontact 579 1083 583 1089 1 vdd
rlabel polycontact 394 1032 398 1036 1 CC0
rlabel polycontact 394 1077 398 1081 1 CC0
rlabel pdcontact 405 1070 409 1074 1 CI0
rlabel pdcontact 405 1060 409 1064 1 CI0
rlabel pdcontact 405 1052 409 1056 1 CI1
rlabel ndcontact 405 1033 409 1037 1 CI1
rlabel polycontact 462 1038 466 1042 1 CI1
rlabel ndcontact 475 1018 479 1022 1 CI2
rlabel ndcontact 475 1034 479 1038 1 CI2
rlabel ndcontact 474 1043 478 1047 1 CI3
rlabel pdcontact 474 1074 478 1078 1 CI3
rlabel polycontact 520 1081 524 1085 1 CI3
rlabel polycontact 519 1016 523 1020 1 CI3
rlabel ndcontact 532 1021 536 1025 1 CI4
rlabel ndcontact 532 1037 536 1041 1 CI4
rlabel ndcontact 531 1046 535 1050 1 CI5
rlabel pdcontact 531 1077 535 1081 1 CI5
rlabel polycontact 580 1059 584 1063 1 CI5
rlabel ndcontact 587 1052 591 1056 1 C0
rlabel pdcontact 587 1084 591 1088 1 C0
rlabel m2contact 618 993 623 998 1 A0
rlabel nwell 973 894 975 896 1 vdd
rlabel pdcontact 959 886 963 892 1 vdd
rlabel nwell 973 842 975 844 1 vdd
rlabel pdcontact 959 834 963 840 1 vdd
rlabel nwell 1062 877 1064 879 1 vdd
rlabel pdcontact 1048 869 1052 875 1 vdd
rlabel ndcontact 1048 851 1052 855 1 gnd
rlabel ndcontact 959 868 963 872 1 gnd
rlabel ndcontact 959 816 963 820 1 gnd
rlabel polycontact 959 823 963 827 1 B1
rlabel ndcontact 967 817 971 821 1 B1N1
rlabel pdcontact 967 834 971 840 1 B1N1
rlabel polycontact 960 875 964 879 1 A1
rlabel ndcontact 967 869 971 873 1 A1N1
rlabel pdcontact 967 886 971 892 1 A1N1
rlabel polycontact 1019 830 1023 834 1 B1N1
rlabel ndcontact 1014 839 1018 844 1 A1N1
rlabel polycontact 1019 871 1023 876 1 B1
rlabel ndcontact 1014 880 1018 885 1 A1
rlabel ndcontact 1031 840 1035 844 1 X1
rlabel ndcontact 1031 881 1035 885 1 X1
rlabel polycontact 1049 858 1053 862 1 X1
rlabel pdcontact 1056 869 1060 875 1 P1
rlabel ndcontact 1056 852 1060 856 1 P1
rlabel polycontact 789 829 793 833 1 clk
rlabel polycontact 790 894 794 898 1 clk
rlabel polycontact 846 857 850 861 1 clk
rlabel metal1 790 909 815 913 1 vdd
rlabel metal1 849 912 874 916 5 vdd
rlabel metal1 898 911 923 915 5 vdd
rlabel metal1 843 909 877 913 1 vdd
rlabel metal1 786 907 820 911 1 vdd
rlabel metal1 899 911 924 913 5 vdd
rlabel nwell 865 903 868 906 1 vdd
rlabel nwell 808 900 811 903 1 vdd
rlabel nwell 920 906 923 909 7 vdd
rlabel ndcontact 802 825 806 829 1 gnd
rlabel ndcontact 859 828 863 832 1 gnd
rlabel ndcontact 906 867 910 871 1 gnd
rlabel pdcontact 801 898 805 902 1 vdd
rlabel pdcontact 858 901 862 905 1 vdd
rlabel pdcontact 906 899 910 905 1 vdd
rlabel ndcontact 914 868 918 872 1 A1
rlabel pdcontact 914 900 918 904 1 A1
rlabel polycontact 789 854 793 858 1 QC1
rlabel pdcontact 801 890 805 894 1 QC3
rlabel ndcontact 801 859 805 863 1 QC3
rlabel polycontact 846 832 850 836 1 QC3
rlabel polycontact 847 897 851 901 1 QC3
rlabel ndcontact 802 834 806 838 1 QC4
rlabel ndcontact 802 850 806 854 1 QC4
rlabel ndcontact 859 837 863 841 1 QC5
rlabel ndcontact 859 853 863 857 1 QC5
rlabel ndcontact 858 862 862 866 1 QC6
rlabel pdcontact 858 893 862 897 1 QC6
rlabel polycontact 907 875 911 879 1 QC6
rlabel nwell 1439 1284 1441 1286 1 vdd
rlabel pdcontact 1425 1276 1429 1282 1 vdd
rlabel nwell 1439 1232 1441 1234 1 vdd
rlabel pdcontact 1425 1224 1429 1230 1 vdd
rlabel nwell 1528 1267 1530 1269 1 vdd
rlabel pdcontact 1514 1259 1518 1265 1 vdd
rlabel ndcontact 1514 1241 1518 1245 1 gnd
rlabel ndcontact 1425 1258 1429 1262 1 gnd
rlabel ndcontact 1425 1206 1429 1210 1 gnd
rlabel polycontact 1425 1213 1429 1217 1 B2
rlabel pdcontact 1433 1224 1437 1230 1 B2N1
rlabel ndcontact 1433 1207 1437 1211 1 B2N1
rlabel polycontact 1426 1265 1430 1269 1 A2
rlabel ndcontact 1433 1259 1437 1263 1 A2N1
rlabel pdcontact 1433 1276 1437 1282 1 A2N1
rlabel ndcontact 1480 1229 1484 1235 1 A2N1
rlabel polycontact 1485 1220 1489 1224 1 B2N1
rlabel polycontact 1485 1261 1489 1266 1 B2
rlabel ndcontact 1480 1270 1484 1275 1 A2
rlabel ndcontact 1497 1230 1501 1235 1 X2
rlabel ndcontact 1497 1271 1501 1276 1 X2
rlabel polycontact 1515 1248 1519 1252 1 X2
rlabel ndcontact 1522 1242 1526 1246 1 P2
rlabel pdcontact 1522 1259 1526 1265 1 P2
rlabel m123contact 1551 1245 1555 1249 1 P2
rlabel pdcontact 1586 1135 1590 1147 1 vdd
rlabel ndcontact 1602 1040 1606 1046 1 gnd
rlabel ndcontact 1579 1053 1583 1059 1 gnd
rlabel ndcontact 1631 1068 1635 1072 1 gnd
rlabel pdcontact 1631 1086 1635 1092 1 vdd
rlabel nwell 1645 1094 1647 1096 1 vdd
rlabel nwell 1603 1138 1607 1142 1 vdd
rlabel polycontact 1572 1046 1576 1050 1 G2
rlabel polycontact 1579 1150 1583 1154 1 G2
rlabel polycontact 1595 1033 1599 1037 1 P2
rlabel polycontact 1571 1116 1575 1120 1 P2
rlabel polycontact 1602 1094 1606 1098 1 G1
rlabel polycontact 1595 1075 1599 1079 1 G1
rlabel pdcontact 1578 1104 1582 1108 1 V2
rlabel pdcontact 1578 1138 1582 1142 1 V2
rlabel pdcontact 1601 1104 1605 1108 1 V2
rlabel ndcontact 1594 1067 1598 1071 1 U2
rlabel ndcontact 1594 1041 1598 1045 1 U2
rlabel pdcontact 1570 1104 1574 1110 1 KC
rlabel ndcontact 1571 1053 1575 1059 1 KC
rlabel polycontact 1632 1075 1636 1079 1 KC
rlabel pdcontact 1609 1104 1613 1110 1 KC
rlabel ndcontact 1602 1066 1606 1072 1 KC
rlabel ndcontact 1639 1069 1643 1073 1 KK
rlabel pdcontact 1639 1086 1643 1092 1 KK
rlabel pdcontact 1726 1115 1730 1127 1 vdd
rlabel pdcontact 1745 1133 1749 1145 1 vdd
rlabel pdcontact 1765 1147 1769 1159 1 vdd
rlabel ndcontact 1749 1033 1753 1042 1 gnd
rlabel polycontact 1766 1162 1770 1166 1 P2
rlabel polycontact 1750 1045 1754 1049 1 P2
rlabel polycontact 1727 1130 1731 1134 1 C1
rlabel polycontact 1750 1093 1754 1097 1 C1
rlabel polycontact 1746 1148 1750 1152 1 P1
rlabel polycontact 1750 1054 1754 1058 1 P1
rlabel ndcontact 1757 1064 1761 1068 1 MP
rlabel ndcontact 1757 1036 1761 1040 1 MP
rlabel ndcontact 1749 1062 1753 1066 1 UP
rlabel ndcontact 1749 1083 1753 1087 1 UP
rlabel pdcontact 1734 1118 1738 1122 1 KP
rlabel pdcontact 1753 1138 1757 1142 1 KP
rlabel pdcontact 1773 1151 1777 1155 1 KP
rlabel ndcontact 1757 1083 1761 1087 1 KP
rlabel metal1 1343 1290 1368 1294 5 vdd
rlabel metal1 1344 1290 1369 1292 5 vdd
rlabel nwell 1365 1285 1368 1288 7 vdd
rlabel ndcontact 1351 1246 1355 1250 1 gnd
rlabel pdcontact 1351 1278 1355 1284 1 vdd
rlabel polycontact 1307 1236 1311 1240 1 clk
rlabel metal1 1310 1291 1335 1295 5 vdd
rlabel metal1 1304 1288 1338 1292 1 vdd
rlabel nwell 1326 1282 1329 1285 1 vdd
rlabel ndcontact 1320 1207 1324 1211 1 gnd
rlabel pdcontact 1319 1280 1323 1284 1 vdd
rlabel pdcontact 1273 1277 1277 1281 1 vdd
rlabel ndcontact 1274 1204 1278 1208 1 gnd
rlabel nwell 1280 1279 1283 1282 1 vdd
rlabel metal1 1258 1286 1292 1290 1 vdd
rlabel metal1 1262 1288 1287 1292 1 vdd
rlabel polycontact 1262 1273 1266 1277 1 clk
rlabel polycontact 1261 1208 1265 1212 1 clk
rlabel polycontact 1221 1254 1225 1258 1 clk
rlabel metal1 1216 1283 1252 1287 5 vdd
rlabel metal1 1216 1283 1252 1286 1 vdd
rlabel nwell 1246 1278 1249 1281 1 vdd
rlabel pdcontact 1232 1273 1236 1277 1 vdd
rlabel ndcontact 1232 1220 1236 1224 1 gnd
rlabel ndcontact 1359 1247 1363 1251 1 A2
rlabel pdcontact 1359 1279 1363 1283 1 A2
rlabel polycontact 1221 1227 1225 1231 1 AA2
rlabel polycontact 1221 1272 1225 1276 1 AA2
rlabel ndcontact 1232 1228 1236 1232 1 R1D
rlabel pdcontact 1232 1247 1236 1251 1 R1D
rlabel polycontact 1261 1233 1265 1237 1 R1D
rlabel pdcontact 1232 1255 1236 1259 1 R2D
rlabel pdcontact 1232 1265 1236 1269 1 R2D
rlabel ndcontact 1274 1213 1278 1217 1 R3D
rlabel ndcontact 1274 1229 1278 1233 1 R3D
rlabel ndcontact 1273 1238 1277 1242 1 R4D
rlabel pdcontact 1273 1269 1277 1273 1 R4D
rlabel polycontact 1308 1276 1312 1280 1 R4D
rlabel polycontact 1307 1211 1311 1215 1 R4D
rlabel ndcontact 1320 1216 1324 1220 1 R5D
rlabel ndcontact 1320 1232 1324 1236 1 R5D
rlabel ndcontact 1319 1241 1323 1245 1 R6D
rlabel pdcontact 1319 1272 1323 1276 1 R6D
rlabel polycontact 1352 1254 1356 1258 1 R6D
rlabel nwell 1134 891 1136 893 1 vdd
rlabel pdcontact 1120 883 1124 889 1 vdd
rlabel nwell 1134 839 1136 841 1 vdd
rlabel pdcontact 1120 831 1124 837 1 vdd
rlabel nwell 1223 874 1225 876 1 vdd
rlabel pdcontact 1209 866 1213 872 1 vdd
rlabel ndcontact 1209 848 1213 852 1 gnd
rlabel ndcontact 1120 865 1124 869 1 gnd
rlabel ndcontact 1120 813 1124 817 1 gnd
rlabel polycontact 1121 872 1125 876 1 P1
rlabel polycontact 1120 820 1124 824 1 C1
rlabel pdcontact 1128 831 1132 837 1 C1N1
rlabel ndcontact 1128 814 1132 818 1 C1N1
rlabel polycontact 1180 827 1184 831 1 C1N1
rlabel ndcontact 1128 866 1132 870 1 P1N1
rlabel pdcontact 1128 883 1132 889 1 P1N1
rlabel ndcontact 1175 836 1179 841 1 P1N1
rlabel polycontact 1180 868 1184 873 1 C1
rlabel ndcontact 1192 837 1196 841 1 S1N
rlabel ndcontact 1192 878 1196 882 1 S1N
rlabel polycontact 1210 855 1214 859 1 S1N
rlabel ndcontact 1217 849 1221 853 1 S1
rlabel pdcontact 1217 866 1221 872 1 S1
rlabel ndcontact 1175 877 1179 883 1 P1
rlabel polycontact 1253 851 1257 855 1 clk
rlabel metal1 1248 880 1284 884 5 vdd
rlabel metal1 1248 880 1284 883 1 vdd
rlabel nwell 1278 875 1281 878 1 vdd
rlabel pdcontact 1264 870 1268 874 1 vdd
rlabel ndcontact 1264 817 1268 821 1 gnd
rlabel polycontact 1253 869 1257 873 1 S1
rlabel polycontact 1253 824 1257 828 1 S1
rlabel ndcontact 1264 825 1268 829 1 TT1
rlabel pdcontact 1264 844 1268 848 1 TT1
rlabel pdcontact 1264 852 1268 856 1 TT2
rlabel pdcontact 1264 862 1268 866 1 TT2
rlabel polycontact 744 875 748 879 1 clk
rlabel metal1 739 904 775 908 5 vdd
rlabel metal1 739 904 775 907 1 vdd
rlabel nwell 769 899 772 902 1 vdd
rlabel pdcontact 755 894 759 898 1 vdd
rlabel ndcontact 755 841 759 845 1 gnd
rlabel polycontact 744 893 748 897 1 AA1
rlabel polycontact 744 848 748 852 1 AA1
rlabel ndcontact 755 849 759 853 1 QC1
rlabel pdcontact 755 868 759 872 1 QC1
rlabel pdcontact 755 876 759 880 1 QC2
rlabel pdcontact 755 886 759 890 1 QC2
rlabel nwell 2121 821 2123 823 1 vdd
rlabel pdcontact 2107 813 2111 819 1 vdd
rlabel nwell 2121 769 2123 771 1 vdd
rlabel pdcontact 2107 761 2111 767 1 vdd
rlabel nwell 2210 804 2212 806 1 vdd
rlabel pdcontact 2196 796 2200 802 1 vdd
rlabel ndcontact 2196 778 2200 782 1 gnd
rlabel ndcontact 2107 795 2111 799 1 gnd
rlabel ndcontact 2107 743 2111 747 1 gnd
rlabel nwell 1861 824 1863 826 1 vdd
rlabel pdcontact 1847 816 1851 822 1 vdd
rlabel nwell 1861 772 1863 774 1 vdd
rlabel pdcontact 1847 764 1851 770 1 vdd
rlabel nwell 1950 807 1952 809 1 vdd
rlabel pdcontact 1936 799 1940 805 1 vdd
rlabel ndcontact 1936 781 1940 785 1 gnd
rlabel ndcontact 1847 798 1851 802 1 gnd
rlabel ndcontact 1847 746 1851 750 1 gnd
rlabel nwell 1880 631 1884 635 1 vdd
rlabel ndcontact 1868 553 1872 559 1 gnd
rlabel pdcontact 1852 628 1856 634 1 vdd
rlabel pdcontact 1878 612 1882 618 1 vdd
rlabel polycontact 1847 753 1851 757 1 B3
rlabel m2contact 1836 588 1840 592 1 B3
rlabel polycontact 1861 588 1865 592 1 B3
rlabel polycontact 1853 621 1857 625 1 B3
rlabel polycontact 1907 801 1911 806 1 B3
rlabel polycontact 1848 805 1852 809 1 A3
rlabel ndcontact 1902 810 1906 815 1 A3
rlabel polycontact 1879 621 1883 625 1 A3
rlabel polycontact 1861 546 1865 550 1 A3
rlabel pdcontact 1860 629 1864 633 1 M4
rlabel ndcontact 1868 580 1872 584 1 M4
rlabel pdcontact 1886 612 1890 616 1 M4
rlabel ndcontact 1860 580 1864 584 1 K4
rlabel ndcontact 1860 554 1864 558 1 K4
rlabel pdcontact 1855 764 1859 770 1 B3N1
rlabel ndcontact 1855 747 1859 751 1 B3N1
rlabel polycontact 1907 760 1911 764 1 B3N1
rlabel ndcontact 1855 799 1859 803 1 A3N1
rlabel pdcontact 1855 816 1859 822 1 A3N1
rlabel ndcontact 1902 769 1906 775 1 A3N1
rlabel ndcontact 1919 769 1923 775 1 X3
rlabel ndcontact 1919 810 1923 816 1 X3
rlabel polycontact 1937 788 1941 792 1 X3
rlabel ndcontact 1944 782 1948 786 1 P3
rlabel pdcontact 1944 799 1948 805 1 P3
rlabel polycontact 2108 802 2112 806 1 P3
rlabel ndcontact 2115 796 2119 800 1 P3N1
rlabel pdcontact 2115 813 2119 819 1 P3N1
rlabel ndcontact 2162 766 2166 772 1 P3N1
rlabel polycontact 2107 750 2111 754 1 C3
rlabel pdcontact 2115 761 2119 767 1 C3N1
rlabel ndcontact 2115 744 2119 748 1 C3N1
rlabel polycontact 2167 757 2171 761 1 C3N1
rlabel polycontact 2167 798 2171 803 1 C3
rlabel ndcontact 2162 807 2166 813 1 P3
rlabel ndcontact 2179 767 2183 772 1 S3N
rlabel ndcontact 2179 808 2183 813 1 S3N
rlabel polycontact 2197 785 2201 789 1 S3N
rlabel ndcontact 2204 779 2208 783 1 S3
rlabel pdcontact 2204 796 2208 802 1 S3
rlabel pdcontact 2030 629 2034 641 1 vdd
rlabel pdcontact 2049 647 2053 659 1 vdd
rlabel pdcontact 2069 661 2073 673 1 vdd
rlabel polycontact 2054 568 2058 572 1 P2
rlabel polycontact 2050 662 2054 666 1 P2
rlabel pdcontact 2086 681 2090 693 1 vdd
rlabel polycontact 2087 696 2091 700 1 P3
rlabel polycontact 2070 676 2074 680 1 P1
rlabel polycontact 2054 559 2058 563 1 P1
rlabel polycontact 2054 520 2058 524 1 P3
rlabel polycontact 2031 644 2035 648 1 C1
rlabel polycontact 2054 607 2058 611 1 C1
rlabel pdcontact 2094 684 2098 690 1 AF
rlabel pdcontact 2077 664 2081 670 1 AF
rlabel pdcontact 2057 651 2061 657 1 AF
rlabel pdcontact 2038 631 2042 637 1 AF
rlabel ndcontact 2061 596 2065 602 1 AF
rlabel ndcontact 2053 596 2057 602 1 LO
rlabel ndcontact 2053 575 2057 581 1 LO
rlabel ndcontact 2061 577 2065 583 1 VE
rlabel ndcontact 2061 549 2065 555 1 VE
rlabel ndcontact 2053 549 2057 555 1 GA
rlabel ndcontact 2053 528 2057 534 1 GA
rlabel ndcontact 2061 530 2065 536 1 gnd
rlabel pdcontact 2195 657 2199 669 1 vdd
rlabel ndcontact 2211 562 2215 568 1 gnd
rlabel ndcontact 2188 575 2192 581 1 gnd
rlabel ndcontact 2240 590 2244 594 1 gnd
rlabel pdcontact 2240 608 2244 614 1 vdd
rlabel nwell 2254 616 2256 618 1 vdd
rlabel nwell 2212 660 2216 664 1 vdd
rlabel pdcontact 2440 658 2444 670 1 vdd
rlabel ndcontact 2458 602 2462 606 1 gnd
rlabel ndcontact 2432 596 2436 600 1 gnd
rlabel polycontact 2188 672 2192 676 1 G3
rlabel pdcontact 2187 660 2191 664 1 V3
rlabel pdcontact 2187 626 2191 630 1 V3
rlabel pdcontact 2210 626 2214 630 1 V3
rlabel polycontact 2180 638 2184 642 1 P3
rlabel polycontact 2204 555 2208 559 1 P3
rlabel polycontact 2211 616 2215 620 1 G2
rlabel polycontact 2204 597 2208 601 1 G2
rlabel ndcontact 2203 589 2207 593 1 U3
rlabel ndcontact 2203 563 2207 567 1 U3
rlabel ndcontact 2180 575 2184 581 1 KJ
rlabel pdcontact 2179 626 2183 632 1 KJ
rlabel pdcontact 2218 626 2222 632 1 KJ
rlabel ndcontact 2211 588 2215 594 1 KJ
rlabel polycontact 2241 597 2245 601 1 KJ
rlabel ndcontact 2248 591 2252 595 1 HQ
rlabel pdcontact 2248 608 2252 614 1 HQ
rlabel m123contact 2415 603 2420 608 1 HQ
rlabel polycontact 2433 604 2437 608 1 HQ
rlabel m123contact 2415 641 2419 645 1 HQ
rlabel polycontact 2441 641 2445 645 1 HQ
rlabel pdcontact 2448 661 2452 667 1 I2
rlabel pdcontact 2448 630 2452 636 1 I2
rlabel pdcontact 2440 628 2444 634 1 OJ
rlabel ndcontact 2440 595 2444 601 1 OJ
rlabel ndcontact 2450 602 2454 608 1 OJ
rlabel metal1 1788 841 1813 845 5 vdd
rlabel metal1 1789 841 1814 843 5 vdd
rlabel nwell 1810 836 1813 839 7 vdd
rlabel ndcontact 1796 797 1800 801 1 gnd
rlabel pdcontact 1796 829 1800 835 1 vdd
rlabel polycontact 1752 787 1756 791 1 clk
rlabel metal1 1755 842 1780 846 5 vdd
rlabel metal1 1749 839 1783 843 1 vdd
rlabel nwell 1771 833 1774 836 1 vdd
rlabel ndcontact 1765 758 1769 762 1 gnd
rlabel pdcontact 1764 831 1768 835 1 vdd
rlabel pdcontact 1718 828 1722 832 1 vdd
rlabel ndcontact 1719 755 1723 759 1 gnd
rlabel nwell 1725 830 1728 833 1 vdd
rlabel metal1 1703 837 1737 841 1 vdd
rlabel metal1 1707 839 1732 843 1 vdd
rlabel polycontact 1707 824 1711 828 1 clk
rlabel polycontact 1706 759 1710 763 1 clk
rlabel polycontact 1666 805 1670 809 1 clk
rlabel metal1 1661 834 1697 838 5 vdd
rlabel metal1 1661 834 1697 837 1 vdd
rlabel nwell 1691 829 1694 832 1 vdd
rlabel pdcontact 1677 824 1681 828 1 vdd
rlabel ndcontact 1677 771 1681 775 1 gnd
rlabel metal1 1788 699 1813 703 5 vdd
rlabel metal1 1789 699 1814 701 5 vdd
rlabel nwell 1810 694 1813 697 7 vdd
rlabel ndcontact 1796 655 1800 659 1 gnd
rlabel pdcontact 1796 687 1800 693 1 vdd
rlabel polycontact 1752 645 1756 649 1 clk
rlabel metal1 1755 700 1780 704 5 vdd
rlabel metal1 1749 697 1783 701 1 vdd
rlabel nwell 1771 691 1774 694 1 vdd
rlabel ndcontact 1765 616 1769 620 1 gnd
rlabel pdcontact 1764 689 1768 693 1 vdd
rlabel pdcontact 1718 686 1722 690 1 vdd
rlabel ndcontact 1719 613 1723 617 1 gnd
rlabel nwell 1725 688 1728 691 1 vdd
rlabel metal1 1703 695 1737 699 1 vdd
rlabel metal1 1707 697 1732 701 1 vdd
rlabel polycontact 1707 682 1711 686 1 clk
rlabel polycontact 1706 617 1710 621 1 clk
rlabel polycontact 1666 663 1670 667 1 clk
rlabel metal1 1661 692 1697 696 5 vdd
rlabel metal1 1661 692 1697 695 1 vdd
rlabel nwell 1691 687 1694 690 1 vdd
rlabel pdcontact 1677 682 1681 686 1 vdd
rlabel ndcontact 1677 629 1681 633 1 gnd
rlabel metal1 2352 821 2377 825 5 vdd
rlabel metal1 2353 821 2378 823 5 vdd
rlabel nwell 2374 816 2377 819 7 vdd
rlabel ndcontact 2360 777 2364 781 1 gnd
rlabel pdcontact 2360 809 2364 815 1 vdd
rlabel polycontact 2316 767 2320 771 1 clk
rlabel metal1 2319 822 2344 826 5 vdd
rlabel metal1 2313 819 2347 823 1 vdd
rlabel nwell 2335 813 2338 816 1 vdd
rlabel ndcontact 2329 738 2333 742 1 gnd
rlabel pdcontact 2328 811 2332 815 1 vdd
rlabel pdcontact 2282 808 2286 812 1 vdd
rlabel ndcontact 2283 735 2287 739 1 gnd
rlabel nwell 2289 810 2292 813 1 vdd
rlabel metal1 2267 817 2301 821 1 vdd
rlabel metal1 2271 819 2296 823 1 vdd
rlabel polycontact 2271 804 2275 808 1 clk
rlabel polycontact 2270 739 2274 743 1 clk
rlabel polycontact 2230 785 2234 789 1 clk
rlabel metal1 2225 814 2261 818 5 vdd
rlabel metal1 2225 814 2261 817 1 vdd
rlabel nwell 2255 809 2258 812 1 vdd
rlabel pdcontact 2241 804 2245 808 1 vdd
rlabel ndcontact 2241 751 2245 755 1 gnd
rlabel ndcontact 1804 798 1808 802 1 A3
rlabel pdcontact 1804 830 1808 834 1 A3
rlabel polycontact 1666 823 1670 827 1 AA3
rlabel polycontact 1666 778 1670 782 1 AA3
rlabel ndcontact 1677 779 1681 783 1 OO8
rlabel pdcontact 1677 798 1681 802 1 OO8
rlabel polycontact 1706 784 1710 788 1 OO8
rlabel pdcontact 1677 806 1681 810 1 O18
rlabel pdcontact 1677 816 1681 820 1 O18
rlabel ndcontact 1718 789 1722 793 1 O13
rlabel pdcontact 1718 820 1722 824 1 O13
rlabel polycontact 1753 827 1757 831 1 O13
rlabel polycontact 1752 762 1756 766 1 O13
rlabel ndcontact 1719 764 1723 768 1 O17
rlabel ndcontact 1719 780 1723 784 1 O17
rlabel ndcontact 1765 767 1769 771 1 O27
rlabel ndcontact 1765 783 1769 787 1 O27
rlabel ndcontact 1764 792 1768 796 1 O37
rlabel pdcontact 1764 823 1768 827 1 O37
rlabel polycontact 1797 805 1801 809 1 O37
rlabel ndcontact 1804 656 1808 660 1 B3
rlabel pdcontact 1804 688 1808 692 1 B3
rlabel polycontact 1666 636 1670 640 1 BB3
rlabel polycontact 1666 681 1670 685 1 BB3
rlabel pdcontact 1677 656 1681 660 1 B51
rlabel ndcontact 1677 637 1681 641 1 B51
rlabel polycontact 1706 642 1710 646 1 B51
rlabel pdcontact 1677 664 1681 668 1 B52
rlabel pdcontact 1677 674 1681 678 1 B52
rlabel pdcontact 1718 678 1722 682 1 B53
rlabel ndcontact 1718 647 1722 651 1 B53
rlabel polycontact 1752 620 1756 624 1 B53
rlabel polycontact 1753 685 1757 689 1 B53
rlabel ndcontact 1719 622 1723 626 1 B54
rlabel ndcontact 1719 638 1723 642 1 B54
rlabel ndcontact 1765 625 1769 629 1 B55
rlabel ndcontact 1765 641 1769 645 1 B55
rlabel ndcontact 1764 650 1768 654 1 B56
rlabel pdcontact 1764 681 1768 685 1 B56
rlabel polycontact 1797 663 1801 667 1 B56
rlabel polycontact 2230 758 2234 762 1 S3
rlabel polycontact 2230 803 2234 807 1 S3
rlabel pdcontact 2241 786 2245 790 1 S3L
rlabel pdcontact 2241 796 2245 800 1 S3L
rlabel pdcontact 2241 778 2245 782 1 S4L
rlabel ndcontact 2241 759 2245 763 1 S4L
rlabel polycontact 2270 764 2274 768 1 S4L
rlabel ndcontact 2283 744 2287 748 1 S5L
rlabel ndcontact 2283 760 2287 764 1 S5L
rlabel ndcontact 2282 769 2286 773 1 S6L
rlabel pdcontact 2282 800 2286 804 1 S6L
rlabel polycontact 2317 807 2321 811 1 S6L
rlabel polycontact 2316 742 2320 746 1 S6L
rlabel ndcontact 2329 747 2333 751 1 S7L
rlabel ndcontact 2329 763 2333 767 1 S7L
rlabel ndcontact 2328 772 2332 776 1 S8L
rlabel pdcontact 2328 803 2332 807 1 S8L
rlabel polycontact 2361 785 2365 789 1 S8L
rlabel ndcontact 2368 778 2372 782 1 SS3
rlabel pdcontact 2368 810 2372 814 1 SS3
rlabel ndcontact 1901 562 1905 566 1 gnd
rlabel pdcontact 1901 580 1905 586 1 vdd
rlabel nwell 1915 588 1917 590 1 vdd
rlabel polycontact 1902 569 1906 573 1 M4
rlabel ndcontact 1909 563 1913 567 1 G3
rlabel pdcontact 1909 580 1913 586 1 G3
rlabel ndcontact 1475 1081 1479 1085 1 gnd
rlabel pdcontact 1475 1099 1479 1105 1 vdd
rlabel nwell 1489 1107 1491 1109 1 vdd
rlabel nwell 1458 1150 1462 1154 1 vdd
rlabel ndcontact 1446 1072 1450 1078 1 gnd
rlabel pdcontact 1430 1147 1434 1153 1 vdd
rlabel pdcontact 1456 1131 1460 1137 1 vdd
rlabel m2contact 1414 1107 1418 1111 1 B2
rlabel polycontact 1439 1107 1443 1111 1 B2
rlabel polycontact 1431 1140 1435 1144 1 B2
rlabel polycontact 1439 1065 1443 1069 1 A2
rlabel polycontact 1457 1140 1461 1144 1 A2
rlabel pdcontact 1438 1148 1442 1152 1 M3
rlabel ndcontact 1446 1099 1450 1103 1 M3
rlabel pdcontact 1464 1131 1468 1135 1 M3
rlabel polycontact 1476 1088 1480 1092 1 M3
rlabel ndcontact 1438 1099 1442 1103 1 K3
rlabel ndcontact 1438 1073 1442 1077 1 K3
rlabel ndcontact 1483 1082 1487 1086 1 G2
rlabel pdcontact 1483 1099 1487 1105 1 G2
rlabel metal1 1366 1182 1391 1186 5 vdd
rlabel metal1 1367 1182 1392 1184 5 vdd
rlabel nwell 1388 1177 1391 1180 7 vdd
rlabel ndcontact 1374 1138 1378 1142 1 gnd
rlabel pdcontact 1374 1170 1378 1176 1 vdd
rlabel polycontact 1330 1128 1334 1132 1 clk
rlabel metal1 1333 1183 1358 1187 5 vdd
rlabel metal1 1327 1180 1361 1184 1 vdd
rlabel nwell 1349 1174 1352 1177 1 vdd
rlabel ndcontact 1343 1099 1347 1103 1 gnd
rlabel pdcontact 1342 1172 1346 1176 1 vdd
rlabel pdcontact 1296 1169 1300 1173 1 vdd
rlabel ndcontact 1297 1096 1301 1100 1 gnd
rlabel nwell 1303 1171 1306 1174 1 vdd
rlabel metal1 1281 1178 1315 1182 1 vdd
rlabel metal1 1285 1180 1310 1184 1 vdd
rlabel polycontact 1285 1165 1289 1169 1 clk
rlabel polycontact 1284 1100 1288 1104 1 clk
rlabel polycontact 1244 1146 1248 1150 1 clk
rlabel metal1 1239 1175 1275 1179 5 vdd
rlabel metal1 1239 1175 1275 1178 1 vdd
rlabel nwell 1269 1170 1272 1173 1 vdd
rlabel pdcontact 1255 1165 1259 1169 1 vdd
rlabel ndcontact 1255 1112 1259 1116 1 gnd
rlabel pdcontact 1382 1171 1386 1175 1 B2
rlabel ndcontact 1382 1139 1386 1143 1 B2
rlabel polycontact 1244 1164 1248 1168 1 BB2
rlabel polycontact 1244 1119 1248 1123 1 BB2
rlabel ndcontact 1255 1120 1259 1124 1 G1A
rlabel pdcontact 1255 1139 1259 1143 1 G1A
rlabel polycontact 1284 1125 1288 1129 1 G1A
rlabel pdcontact 1255 1147 1259 1151 1 G2A
rlabel pdcontact 1255 1157 1259 1161 1 G2A
rlabel ndcontact 1297 1105 1301 1109 1 G3A
rlabel ndcontact 1297 1121 1301 1125 1 G3A
rlabel ndcontact 1296 1130 1300 1134 1 G4A
rlabel pdcontact 1296 1161 1300 1165 1 G4A
rlabel polycontact 1331 1168 1335 1172 1 G4A
rlabel polycontact 1330 1103 1334 1107 1 G4A
rlabel ndcontact 1343 1108 1347 1112 1 G5A
rlabel ndcontact 1343 1124 1347 1128 1 G5A
rlabel ndcontact 1342 1133 1346 1137 1 G6A
rlabel pdcontact 1342 1164 1346 1168 1 G6A
rlabel polycontact 1375 1146 1379 1150 1 G6A
rlabel m3contact 2160 719 2165 724 1 P3
rlabel pdcontact 2569 658 2573 670 1 vdd
rlabel ndcontact 2587 602 2591 606 1 gnd
rlabel ndcontact 2561 596 2565 600 1 gnd
rlabel pdcontact 2577 661 2581 667 1 I3
rlabel pdcontact 2577 630 2581 636 1 I3
rlabel metal1 2767 677 2792 681 5 vdd
rlabel metal1 2768 677 2793 679 5 vdd
rlabel nwell 2789 672 2792 675 7 vdd
rlabel ndcontact 2775 633 2779 637 1 gnd
rlabel pdcontact 2775 665 2779 671 1 vdd
rlabel polycontact 2731 623 2735 627 1 clk
rlabel metal1 2734 678 2759 682 5 vdd
rlabel metal1 2728 675 2762 679 1 vdd
rlabel nwell 2750 669 2753 672 1 vdd
rlabel ndcontact 2744 594 2748 598 1 gnd
rlabel pdcontact 2743 667 2747 671 1 vdd
rlabel pdcontact 2697 664 2701 668 1 vdd
rlabel ndcontact 2698 591 2702 595 1 gnd
rlabel nwell 2704 666 2707 669 1 vdd
rlabel metal1 2682 673 2716 677 1 vdd
rlabel metal1 2686 675 2711 679 1 vdd
rlabel polycontact 2686 660 2690 664 1 clk
rlabel polycontact 2685 595 2689 599 1 clk
rlabel polycontact 2645 641 2649 645 1 clk
rlabel metal1 2640 670 2676 674 5 vdd
rlabel metal1 2640 670 2676 673 1 vdd
rlabel nwell 2670 665 2673 668 1 vdd
rlabel pdcontact 2656 660 2660 664 1 vdd
rlabel ndcontact 2656 607 2660 611 1 gnd
rlabel polycontact 2645 614 2649 618 1 C4
rlabel polycontact 2645 659 2649 663 1 C4
rlabel pdcontact 2656 652 2660 656 1 9R
rlabel pdcontact 2656 642 2660 646 1 9R
rlabel pdcontact 2656 634 2660 638 1 9W
rlabel ndcontact 2656 615 2660 619 1 9W
rlabel polycontact 2685 620 2689 624 1 9W
rlabel ndcontact 2698 600 2702 604 1 9T
rlabel ndcontact 2698 616 2702 620 1 9T
rlabel ndcontact 2697 625 2701 629 1 9P
rlabel pdcontact 2697 656 2701 660 1 9P
rlabel polycontact 2731 598 2735 602 1 9P
rlabel polycontact 2732 663 2736 667 1 9P
rlabel ndcontact 2744 603 2748 607 1 9E
rlabel ndcontact 2744 619 2748 623 1 9E
rlabel ndcontact 2743 628 2747 632 1 9V
rlabel pdcontact 2743 659 2747 663 1 9V
rlabel polycontact 2776 641 2780 645 1 9V
rlabel ndcontact 2783 634 2787 638 1 CC4
rlabel pdcontact 2783 666 2787 670 1 CC4
rlabel ndcontact 2603 607 2607 611 1 gnd
rlabel pdcontact 2603 625 2607 631 1 vdd
rlabel nwell 2617 633 2619 635 1 vdd
rlabel ndcontact 2569 595 2573 601 1 C4N
rlabel ndcontact 2579 602 2583 608 1 C4N
rlabel pdcontact 2569 628 2573 634 1 C4N
rlabel polycontact 2604 614 2608 618 1 C4N
rlabel ndcontact 2611 608 2615 612 1 C4
rlabel pdcontact 2611 625 2615 631 1 C4
rlabel ndcontact 2485 607 2489 611 1 gnd
rlabel pdcontact 2485 625 2489 631 1 vdd
rlabel nwell 2499 633 2501 635 1 vdd
rlabel polycontact 2486 614 2490 618 1 OJ
rlabel ndcontact 2493 608 2497 612 1 ZC
rlabel pdcontact 2493 625 2497 631 1 ZC
rlabel m2contact 2525 605 2529 607 1 ZC
rlabel polycontact 2562 604 2566 608 1 ZC
rlabel polycontact 2570 673 2574 677 1 ZC
rlabel pdcontact 1868 1136 1872 1148 1 vdd
rlabel ndcontact 1886 1080 1890 1084 1 gnd
rlabel ndcontact 1860 1074 1864 1078 1 gnd
rlabel pdcontact 1876 1108 1880 1114 1 I0
rlabel pdcontact 1876 1139 1880 1145 1 I0
rlabel m123contact 1844 1082 1846 1085 1 KK
rlabel m123contact 1844 1119 1846 1122 1 KK
rlabel polycontact 1869 1119 1873 1123 1 KK
rlabel polycontact 1861 1082 1865 1086 1 KK
rlabel nwell 1915 1123 1917 1125 1 vdd
rlabel pdcontact 1901 1115 1905 1121 1 vdd
rlabel ndcontact 1901 1097 1905 1101 1 gnd
rlabel ndcontact 1878 1080 1882 1086 1 C3N
rlabel ndcontact 1868 1073 1872 1079 1 C3N
rlabel pdcontact 1868 1106 1872 1112 1 C3N
rlabel polycontact 1902 1104 1906 1108 1 C3N
rlabel pdcontact 1909 1115 1913 1121 1 C3
rlabel ndcontact 1909 1098 1913 1102 1 C3
rlabel nwell 1819 1120 1821 1122 1 vdd
rlabel pdcontact 1805 1112 1809 1118 1 vdd
rlabel ndcontact 1805 1094 1809 1098 1 gnd
rlabel polycontact 1806 1101 1810 1105 1 KP
rlabel pdcontact 1813 1112 1817 1118 1 PP
rlabel ndcontact 1813 1095 1817 1099 1 PP
rlabel polycontact 1869 1151 1873 1155 1 PP
rlabel polycontact 1879 1073 1883 1077 1 PP
rlabel pdcontact 2306 637 2310 649 1 vdd
rlabel pdcontact 2325 655 2329 667 1 vdd
rlabel pdcontact 2345 669 2349 681 1 vdd
rlabel ndcontact 2329 555 2333 564 1 gnd
rlabel polycontact 2346 684 2350 688 1 P3
rlabel polycontact 2330 567 2334 571 1 P3
rlabel polycontact 2330 576 2334 580 1 P2
rlabel polycontact 2326 670 2330 674 1 P2
rlabel polycontact 2307 652 2311 656 1 G1
rlabel polycontact 2330 615 2334 619 1 G1
rlabel ndcontact 2337 558 2341 562 1 AW
rlabel ndcontact 2337 586 2341 590 1 AW
rlabel ndcontact 2329 584 2333 588 1 NT
rlabel ndcontact 2329 605 2333 609 1 NT
rlabel ndcontact 2337 605 2341 609 1 LT
rlabel pdcontact 2314 640 2318 644 1 LT
rlabel pdcontact 2333 660 2337 664 1 LT
rlabel pdcontact 2353 673 2357 677 1 LT
rlabel ndcontact 2381 616 2385 620 1 gnd
rlabel pdcontact 2381 634 2385 640 1 vdd
rlabel nwell 2395 642 2397 644 1 vdd
rlabel polycontact 2382 623 2386 627 1 LT
rlabel ndcontact 2389 617 2393 621 1 LTT
rlabel pdcontact 2389 634 2393 640 1 LTT
rlabel polycontact 2451 595 2455 599 1 LTT
rlabel polycontact 2441 673 2445 677 1 LTT
rlabel nwell 2127 530 2129 532 1 vdd
rlabel pdcontact 2113 522 2117 528 1 vdd
rlabel ndcontact 2113 504 2117 508 1 gnd
rlabel polycontact 2114 511 2118 515 1 AF
rlabel pdcontact 2121 522 2125 528 1 HE
rlabel ndcontact 2121 505 2125 509 1 HE
rlabel polycontact 2580 595 2584 599 1 HE
rlabel polycontact 2570 641 2574 645 1 HE
rlabel polycontact 2181 568 2185 572 1 G3
rlabel nwell 1630 1281 1632 1283 1 vdd
rlabel pdcontact 1616 1273 1620 1279 1 vdd
rlabel nwell 1630 1229 1632 1231 1 vdd
rlabel pdcontact 1616 1221 1620 1227 1 vdd
rlabel nwell 1719 1264 1721 1266 1 vdd
rlabel pdcontact 1705 1256 1709 1262 1 vdd
rlabel ndcontact 1705 1238 1709 1242 1 gnd
rlabel ndcontact 1616 1255 1620 1259 1 gnd
rlabel ndcontact 1616 1203 1620 1207 1 gnd
rlabel polycontact 1617 1262 1621 1266 1 P2
rlabel ndcontact 1624 1256 1628 1260 1 P2N1
rlabel pdcontact 1624 1273 1628 1279 1 P2N1
rlabel ndcontact 1671 1226 1675 1232 1 P2N1
rlabel polycontact 1616 1210 1620 1214 1 C2
rlabel pdcontact 1624 1221 1628 1227 1 C2N1
rlabel ndcontact 1624 1204 1628 1208 1 C2N1
rlabel polycontact 1676 1217 1680 1221 1 C2N1
rlabel polycontact 1676 1258 1680 1263 1 C2
rlabel ndcontact 1688 1227 1692 1232 1 S2N
rlabel ndcontact 1688 1268 1692 1273 1 S2N
rlabel polycontact 1706 1245 1710 1249 1 S2N
rlabel pdcontact 1713 1256 1717 1262 1 S2
rlabel ndcontact 1713 1239 1717 1243 1 S2
rlabel metal1 1861 1291 1886 1295 5 vdd
rlabel metal1 1862 1291 1887 1293 5 vdd
rlabel nwell 1883 1286 1886 1289 7 vdd
rlabel ndcontact 1869 1247 1873 1251 1 gnd
rlabel pdcontact 1869 1279 1873 1285 1 vdd
rlabel polycontact 1825 1237 1829 1241 1 clk
rlabel metal1 1828 1292 1853 1296 5 vdd
rlabel metal1 1822 1289 1856 1293 1 vdd
rlabel nwell 1844 1283 1847 1286 1 vdd
rlabel ndcontact 1838 1208 1842 1212 1 gnd
rlabel pdcontact 1837 1281 1841 1285 1 vdd
rlabel pdcontact 1791 1278 1795 1282 1 vdd
rlabel ndcontact 1792 1205 1796 1209 1 gnd
rlabel nwell 1798 1280 1801 1283 1 vdd
rlabel metal1 1776 1287 1810 1291 1 vdd
rlabel metal1 1780 1289 1805 1293 1 vdd
rlabel polycontact 1780 1274 1784 1278 1 clk
rlabel polycontact 1779 1209 1783 1213 1 clk
rlabel polycontact 1739 1255 1743 1259 1 clk
rlabel metal1 1734 1284 1770 1288 5 vdd
rlabel metal1 1734 1284 1770 1287 1 vdd
rlabel nwell 1764 1279 1767 1282 1 vdd
rlabel pdcontact 1750 1274 1754 1278 1 vdd
rlabel ndcontact 1750 1221 1754 1225 1 gnd
rlabel polycontact 1739 1228 1743 1232 1 S2
rlabel polycontact 1739 1273 1743 1277 1 S2
rlabel pdcontact 1750 1266 1754 1270 1 SK2
rlabel pdcontact 1750 1256 1754 1260 1 SK2
rlabel pdcontact 1750 1248 1754 1252 1 SK3
rlabel ndcontact 1750 1229 1754 1233 1 SK3
rlabel polycontact 1779 1234 1783 1238 1 SK3
rlabel ndcontact 1792 1214 1796 1218 1 SK4
rlabel ndcontact 1792 1230 1796 1234 1 SK4
rlabel ndcontact 1791 1239 1795 1243 1 SK5
rlabel pdcontact 1791 1270 1795 1274 1 SK5
rlabel polycontact 1826 1277 1830 1281 1 SK5
rlabel polycontact 1825 1212 1829 1216 1 SK5
rlabel ndcontact 1838 1217 1842 1221 1 SK6
rlabel ndcontact 1838 1233 1842 1237 1 SK6
rlabel ndcontact 1837 1242 1841 1246 1 SK7
rlabel pdcontact 1837 1273 1841 1277 1 SK7
rlabel polycontact 1870 1255 1874 1259 1 SK7
rlabel ndcontact 1877 1248 1881 1252 1 SS2
rlabel pdcontact 1877 1280 1881 1284 1 SS2
rlabel nwell 758 1261 760 1263 1 vdd
rlabel pdcontact 744 1253 748 1259 1 vdd
rlabel nwell 758 1209 760 1211 1 vdd
rlabel pdcontact 744 1201 748 1207 1 vdd
rlabel nwell 847 1244 849 1246 1 vdd
rlabel pdcontact 833 1236 837 1242 1 vdd
rlabel ndcontact 833 1218 837 1222 1 gnd
rlabel ndcontact 744 1235 748 1239 1 gnd
rlabel ndcontact 744 1183 748 1187 1 gnd
rlabel polycontact 745 1242 749 1246 1 P0
rlabel polycontact 744 1190 748 1194 1 C0
rlabel polycontact 804 1238 808 1243 1 C0
rlabel ndcontact 752 1236 756 1240 1 P0N1
rlabel ndcontact 799 1206 803 1211 1 P0N1
rlabel pdcontact 752 1201 756 1207 1 C0N1
rlabel ndcontact 752 1184 756 1188 1 C0N1
rlabel polycontact 804 1197 808 1201 1 C0N1
rlabel ndcontact 799 1247 803 1252 1 P0
rlabel ndcontact 816 1248 820 1252 1 S0N
rlabel ndcontact 816 1207 820 1211 1 S0N
rlabel polycontact 834 1225 838 1229 1 S0N
rlabel ndcontact 841 1219 845 1223 1 S0
rlabel pdcontact 841 1236 845 1242 1 S0
rlabel pdcontact 752 1253 756 1259 1 P0N1
rlabel polycontact 862 1235 866 1239 1 clk
rlabel polycontact 930 1189 934 1193 1 clk
rlabel polycontact 931 1254 935 1258 1 clk
rlabel polycontact 987 1217 991 1221 1 clk
rlabel metal1 931 1269 956 1273 1 vdd
rlabel metal1 990 1272 1015 1276 5 vdd
rlabel metal1 1039 1271 1064 1275 5 vdd
rlabel metal1 984 1269 1018 1273 1 vdd
rlabel metal1 927 1267 961 1271 1 vdd
rlabel metal1 857 1264 893 1268 5 vdd
rlabel metal1 857 1264 893 1267 1 vdd
rlabel metal1 1040 1271 1065 1273 5 vdd
rlabel nwell 1006 1263 1009 1266 1 vdd
rlabel nwell 949 1260 952 1263 1 vdd
rlabel nwell 887 1259 890 1262 1 vdd
rlabel nwell 1061 1266 1064 1269 7 vdd
rlabel pdcontact 873 1254 877 1258 1 vdd
rlabel ndcontact 873 1201 877 1205 1 gnd
rlabel ndcontact 943 1185 947 1189 1 gnd
rlabel ndcontact 1000 1188 1004 1192 1 gnd
rlabel ndcontact 1047 1227 1051 1231 1 gnd
rlabel pdcontact 942 1258 946 1262 1 vdd
rlabel pdcontact 999 1261 1003 1265 1 vdd
rlabel pdcontact 1047 1259 1051 1265 1 vdd
rlabel polycontact 862 1208 866 1212 1 S0
rlabel polycontact 862 1253 866 1257 1 S0
rlabel pdcontact 873 1246 877 1250 1 SJ0
rlabel pdcontact 873 1236 877 1240 1 SJ0
rlabel pdcontact 873 1228 877 1232 1 SJ1
rlabel ndcontact 873 1209 877 1213 1 SJ1
rlabel polycontact 930 1214 934 1218 1 SJ1
rlabel ndcontact 943 1194 947 1198 1 SJ2
rlabel ndcontact 943 1210 947 1214 1 SJ2
rlabel ndcontact 942 1219 946 1223 1 SJ3
rlabel pdcontact 942 1250 946 1254 1 SJ3
rlabel polycontact 987 1192 991 1196 1 SJ3
rlabel polycontact 988 1257 992 1261 1 SJ3
rlabel ndcontact 1000 1197 1004 1201 1 SJ4
rlabel ndcontact 1000 1213 1004 1217 1 SJ4
rlabel ndcontact 999 1222 1003 1226 1 SJ5
rlabel pdcontact 999 1253 1003 1257 1 SJ5
rlabel polycontact 1048 1235 1052 1239 1 SJ5
rlabel ndcontact 1055 1228 1059 1232 1 SS0
rlabel pdcontact 1055 1260 1059 1264 1 SS0
rlabel polycontact 1297 805 1301 809 1 clk
rlabel polycontact 1298 870 1302 874 1 clk
rlabel polycontact 1354 833 1358 837 1 clk
rlabel metal1 1298 885 1323 889 1 vdd
rlabel metal1 1357 888 1382 892 5 vdd
rlabel metal1 1351 885 1385 889 1 vdd
rlabel metal1 1294 883 1328 887 1 vdd
rlabel nwell 1373 879 1376 882 1 vdd
rlabel nwell 1316 876 1319 879 1 vdd
rlabel ndcontact 1310 801 1314 805 1 gnd
rlabel ndcontact 1367 804 1371 808 1 gnd
rlabel pdcontact 1309 874 1313 878 1 vdd
rlabel pdcontact 1366 877 1370 881 1 vdd
rlabel polycontact 1297 830 1301 834 1 TT1
rlabel ndcontact 1310 810 1314 814 1 TT3
rlabel ndcontact 1310 826 1314 830 1 TT3
rlabel ndcontact 1309 835 1313 839 1 TT4
rlabel pdcontact 1309 866 1313 870 1 TT4
rlabel polycontact 1355 873 1359 877 1 TT4
rlabel polycontact 1354 808 1358 812 1 TT4
rlabel ndcontact 1367 813 1371 817 1 TT5
rlabel ndcontact 1367 829 1371 833 1 TT5
rlabel ndcontact 1366 838 1370 842 1 TT6
rlabel pdcontact 1366 869 1370 873 1 TT6
rlabel metal1 1396 887 1421 891 5 vdd
rlabel metal1 1397 887 1422 889 5 vdd
rlabel nwell 1418 882 1421 885 7 vdd
rlabel ndcontact 1404 843 1408 847 1 gnd
rlabel pdcontact 1404 875 1408 881 1 vdd
rlabel polycontact 1405 851 1409 855 1 TT6
rlabel ndcontact 1412 844 1416 848 1 SS1
rlabel pdcontact 1412 876 1416 880 1 SS1
rlabel pdcontact 990 743 994 749 1 vdd
rlabel pdcontact 964 759 968 765 1 vdd
rlabel ndcontact 980 684 984 690 1 gnd
rlabel nwell 992 762 996 766 1 vdd
rlabel nwell 1023 719 1025 721 1 vdd
rlabel pdcontact 1009 711 1013 717 1 vdd
rlabel ndcontact 1009 693 1013 697 1 gnd
rlabel pdcontact 1120 759 1124 771 1 vdd
rlabel ndcontact 1136 664 1140 670 1 gnd
rlabel ndcontact 1113 677 1117 683 1 gnd
rlabel ndcontact 1165 692 1169 696 1 gnd
rlabel pdcontact 1165 710 1169 716 1 vdd
rlabel nwell 1179 718 1181 720 1 vdd
rlabel pdcontact 1173 710 1177 716 1 C2
rlabel ndcontact 1173 693 1177 697 1 C2
rlabel polycontact 1166 699 1170 703 1 C2N
rlabel ndcontact 1136 690 1140 696 1 C2N
rlabel pdcontact 1143 728 1147 734 1 C2N
rlabel pdcontact 1104 728 1108 734 1 C2N
rlabel ndcontact 1105 677 1109 683 1 C2N
rlabel m2contact 948 719 952 723 1 B1
rlabel polycontact 973 677 977 681 1 A1
rlabel polycontact 991 752 995 756 1 A1
rlabel polycontact 973 719 977 723 1 B1
rlabel polycontact 965 752 969 756 1 B1
rlabel pdcontact 972 760 976 764 1 M2
rlabel ndcontact 980 711 984 715 1 M2
rlabel pdcontact 998 743 1002 747 1 M2
rlabel polycontact 1010 700 1014 704 1 M2
rlabel ndcontact 972 685 976 689 1 K2
rlabel ndcontact 972 711 976 715 1 K2
rlabel pdcontact 1017 711 1021 717 1 G1
rlabel ndcontact 1017 694 1021 698 1 G1
rlabel polycontact 1106 670 1110 674 1 G1
rlabel polycontact 1113 774 1117 778 1 G1
rlabel polycontact 1136 718 1140 722 1 C1
rlabel polycontact 1129 699 1133 703 1 C1
rlabel polycontact 1105 740 1109 744 1 P1
rlabel polycontact 1129 657 1133 661 1 P1
rlabel ndcontact 1128 691 1132 695 1 U1
rlabel ndcontact 1128 665 1132 669 1 U1
rlabel pdcontact 1112 762 1116 766 1 V1
rlabel pdcontact 1112 728 1116 732 1 V1
rlabel pdcontact 1135 728 1139 732 1 V1
rlabel nwell 1137 762 1141 766 1 vdd
rlabel metal1 902 780 927 784 5 vdd
rlabel metal1 903 780 928 782 5 vdd
rlabel nwell 924 775 927 778 7 vdd
rlabel ndcontact 910 736 914 740 1 gnd
rlabel pdcontact 910 768 914 774 1 vdd
rlabel polycontact 863 726 867 730 1 clk
rlabel metal1 866 781 891 785 5 vdd
rlabel metal1 860 778 894 782 1 vdd
rlabel nwell 882 772 885 775 1 vdd
rlabel ndcontact 876 697 880 701 1 gnd
rlabel pdcontact 875 770 879 774 1 vdd
rlabel polycontact 814 698 818 702 1 clk
rlabel polycontact 815 763 819 767 1 clk
rlabel metal1 815 778 840 782 1 vdd
rlabel metal1 811 776 845 780 1 vdd
rlabel nwell 833 769 836 772 1 vdd
rlabel ndcontact 827 694 831 698 1 gnd
rlabel pdcontact 826 767 830 771 1 vdd
rlabel ndcontact 785 710 789 714 1 gnd
rlabel pdcontact 785 763 789 767 1 vdd
rlabel nwell 799 768 802 771 1 vdd
rlabel metal1 769 773 805 776 1 vdd
rlabel metal1 769 773 805 777 5 vdd
rlabel polycontact 774 744 778 748 1 clk
rlabel polycontact 774 762 778 766 1 BB1
rlabel polycontact 774 717 778 721 1 BB1
rlabel pdcontact 785 737 789 741 1 BF1
rlabel ndcontact 785 718 789 722 1 BF1
rlabel polycontact 814 723 818 727 1 BF1
rlabel pdcontact 785 745 789 749 1 BF2
rlabel pdcontact 785 755 789 759 1 BF2
rlabel pdcontact 826 759 830 763 1 BF3
rlabel ndcontact 826 728 830 732 1 BF3
rlabel ndcontact 827 719 831 723 1 BF4
rlabel ndcontact 827 703 831 707 1 BF4
rlabel polycontact 864 766 868 770 1 BF3
rlabel polycontact 863 701 867 705 1 BF3
rlabel ndcontact 876 706 880 710 1 BF5
rlabel ndcontact 876 722 880 726 1 BF5
rlabel ndcontact 875 731 879 735 1 BF6
rlabel pdcontact 875 762 879 766 1 BF6
rlabel polycontact 911 744 915 748 1 BF6
rlabel ndcontact 918 737 922 741 1 B1
rlabel pdcontact 918 769 922 773 1 B1
rlabel m123contact 1084 859 1090 865 1 P1
rlabel ndcontact 1671 1267 1675 1273 1 P2
<< end >>
