* SPICE3 file created from carry.ext - technology: scmos

.option scale=90n

M1000 Z0 P0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1001 P0 X0 gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1002 C2N C1 V1 vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1003 KC G1 V2 vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1004 gnd P2 U2 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1005 I2 HQ OJ vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1006 C4 C4N vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1007 I3 AFF C4N vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1008 B0N1 B0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1009 Z0 C0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1010 KP P2 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1011 AF P3 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1012 C4 C4N gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1013 Z0 C0 M0 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1014 C1 Y0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1015 A0N1 A0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1016 HQ L34 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1017 VE P1 GA Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1018 OJ HQ gnd Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1019 L34 G2 U3 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1020 HQ L34 gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1021 AW P3 gnd Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1022 A0N1 A0 gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1023 C1 Z0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1024 MP P1 UP Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1025 AF C1 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1026 gnd G3 L34 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1027 C2N C1 U1 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1028 AFF AF vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1029 C1 Z0 K0 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1030 gnd P3 GA Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1031 LT P3 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1032 AF C1 LO Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1033 V1 P1 C2N vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1034 I0 KPK vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1035 V2 P2 KC vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1036 Y0 A0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1037 LT G1 NT Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1038 B0N1 B0 gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1039 MP P2 gnd Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1040 gnd B0 N0 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1041 I0 KK C3N vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1042 KK KC vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1043 gnd AFF C4N Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1044 C4N OK gnd Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1045 KP C1 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1046 KC G1 U2 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1047 AF P2 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1048 vdd G3 V3 vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1049 I2 6R vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1050 6R LT vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1051 X0 B0N1 A0N1 Gnd nfet w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1052 gnd 6R OJ Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1053 C2 C2N gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1054 Y0 B0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1055 AF P1 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1056 LT P2 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1057 I3 OK vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1058 gnd P0 M0 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1059 P0 X0 vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1060 vdd G2 V2 vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1061 C3N KK gnd Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1062 LT G1 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1063 L34 G2 V3 vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1064 6R LT gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1065 gnd P3 U3 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1066 gnd G1 C2N Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1067 AFF AF gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1068 X0 B0 A0 Gnd nfet w=6 l=2
+  ad=59.999996p pd=32u as=54p ps=30u
M1069 OK OJ gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1070 gnd P1 U1 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1071 KPK KP vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1072 Y0 A0 N0 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1073 C2 C2N vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1074 KPK KP gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1075 VE P2 LO Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1076 KP P1 vdd vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1077 gnd Y0 K0 Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1078 V3 P3 L34 vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1079 C3 C3N vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1080 AW P2 NT Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1081 C3 C3N gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1082 KK KC gnd Gnd nfet w=3 l=2
+  ad=19p pd=18u as=19p ps=18u
M1083 OK OJ vdd vdd pfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1084 KP C1 UP Gnd nfet w=9 l=2
+  ad=45p pd=28u as=45p ps=28u
M1085 gnd KPK C3N Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
M1086 vdd G1 V1 vdd pfet w=12 l=2
+  ad=59.999996p pd=34u as=59.999996p ps=34u
M1087 gnd G2 KC Gnd nfet w=6 l=2
+  ad=29.999998p pd=22u as=29.999998p ps=22u
C0 G1 P2 0.290858f
C1 U1 m3_937_n361# 2.34e-20
C2 UP MP 0.092785f
C3 Y0 vdd 0.312468f
C4 P3 V3 0.056801f
C5 OK C4N 0.056757f
C6 vdd C4N 0.053819f
C7 C2N m3_937_n361# 2.34e-20
C8 G1 U2 0.041965f
C9 M0 gnd 0.061857f
C10 C3N vdd 0.053754f
C11 P3 AF 7.27e-19
C12 P3 GA 0.055711f
C13 vdd I2 0.149953f
C14 G1 V1 0.055711f
C15 gnd LT 0.056518f
C16 KPK vdd 0.194108f
C17 NT LT 0.092785f
C18 m2_937_n397# m3_937_n361# 0.00709f
C19 vdd V3 0.191129f
C20 I0 KK 0.05668f
C21 C1 K0 0.061857f
C22 C2 vdd 0.094864f
C23 P1 UP 0.055711f
C24 vdd m3_1120_n429# 0.003759f
C25 m2_496_n352# m3_496_n300# 4.06e-19
C26 vdd AF 0.764456f
C27 U3 m3_1717_n374# 2.34e-20
C28 vdd m3_937_n361# 0.003759f
C29 P2 m3_1120_n429# 1.53e-19
C30 U3 P3 0.041965f
C31 HQ AW 3.8e-20
C32 C4N AFF 0.177461f
C33 P2 AF 7.27e-19
C34 C1 P1 0.290858f
C35 AW gnd 0.092785f
C36 KP UP 0.092785f
C37 C0 vdd 0.13033f
C38 U2 m3_1120_n429# 2.34e-20
C39 vdd m2_1123_n465# 0.008839f
C40 NT AW 0.092785f
C41 HQ gnd 0.127318f
C42 vdd m2_1729_n327# 0.008839f
C43 B0 m2_496_n352# 3.61e-19
C44 C3 m3_1503_n436# 1.87e-19
C45 M0 P0 0.055711f
C46 Z0 K0 0.055711f
C47 KP C1 0.264241f
C48 KPK C3N 0.121267f
C49 VE P2 0.05668f
C50 m3_937_n361# V1 1.87e-20
C51 m3_2144_n302# C4 1.87e-19
C52 B0 gnd 0.056518f
C53 U2 m2_1123_n465# 9.6e-20
C54 A0 m2_453_n347# 3.1e-19
C55 G1 m3_937_n361# 0.004826f
C56 AF AFF 0.058778f
C57 U1 C1 0.041965f
C58 MP gnd 0.092785f
C59 A0 vdd 0.405391f
C60 G1 m2_1123_n465# 6.24e-19
C61 LT 6R 0.058778f
C62 LO P2 0.055711f
C63 C2N C1 0.174647f
C64 m3_1717_n374# L34 2.34e-20
C65 KK vdd 0.140896f
C66 K0 gnd 0.061857f
C67 P3 L34 0.041965f
C68 Z0 P0 0.162736f
C69 gnd C4 0.072183f
C70 C3 gnd 0.072183f
C71 KK P2 3.77e-21
C72 C1 m2_937_n397# 6.24e-19
C73 HQ OJ 0.112874f
C74 vdd A0N1 0.094864f
C75 gnd OJ 0.207735f
C76 Y0 N0 0.061857f
C77 KC vdd 0.06532f
C78 P3 LT 7.27e-19
C79 gnd P0 0.072183f
C80 m3_1717_n374# G3 0.002413f
C81 vdd L34 0.06532f
C82 KC P2 0.041965f
C83 Y0 A0 0.11336f
C84 C1 vdd 0.705712f
C85 HQ 6R 0.14318f
C86 OK I3 7.27e-19
C87 m2_1123_n465# m3_1120_n429# 0.00709f
C88 gnd 6R 0.168434f
C89 vdd I3 0.149953f
C90 m2_1729_n327# V3 9.6e-20
C91 KP gnd 0.056518f
C92 KC U2 0.061857f
C93 P1 MP 0.05668f
C94 C1 P2 0.290858f
C95 VE GA 0.092785f
C96 gnd X0 0.080082f
C97 vdd LT 0.518157f
C98 U1 gnd 0.061857f
C99 C3N KK 0.112874f
C100 V2 vdd 0.191129f
C101 KC G1 0.174647f
C102 vdd m3_1503_n436# 0.001729f
C103 AW P3 0.05668f
C104 B0 X0 0.001447f
C105 vdd G3 0.060843f
C106 C1 V1 0.041965f
C107 P2 LT 7.27e-19
C108 KPK KK 0.14318f
C109 V2 P2 0.056801f
C110 C2N gnd 0.118374f
C111 G2 vdd 0.09441f
C112 LO AF 0.092785f
C113 m2_453_n347# m3_496_n300# 0.007496f
C114 vdd m3_2144_n302# 0.001729f
C115 HQ P3 9.58e-19
C116 C1 Y0 0.162736f
C117 P3 gnd 0.054984f
C118 Z0 vdd 0.291414f
C119 B0N1 m2_496_n352# 0.001081f
C120 vdd m3_496_n300# 0.001731f
C121 I3 AFF 0.05668f
C122 G1 LT 0.264241f
C123 U3 m2_1729_n327# 9.6e-20
C124 B0N1 gnd 0.072183f
C125 V2 G1 0.041965f
C126 vdd m2_496_n352# 0.004941f
C127 gnd m2_453_n347# 0.002765f
C128 LO VE 0.092785f
C129 I3 C4N 0.123714f
C130 6R OJ 0.121267f
C131 KP P1 7.27e-19
C132 B0N1 B0 1.62e-19
C133 OK gnd 0.113518f
C134 HQ vdd 0.140896f
C135 AW P2 0.05668f
C136 B0 m2_453_n347# 7.05e-19
C137 KC m3_1120_n429# 2.34e-20
C138 V3 L34 0.247428f
C139 U1 P1 0.041965f
C140 P2 gnd 0.054984f
C141 C3N m3_1503_n436# 1.12e-19
C142 A0 N0 0.055711f
C143 B0 vdd 0.19512f
C144 X0 P0 0.058778f
C145 C1 AF 0.264241f
C146 Z0 Y0 0.227363f
C147 NT P2 0.055711f
C148 C2N P1 0.041965f
C149 m3_2144_n302# C4N 1.12e-19
C150 KC m2_1123_n465# 0.018008f
C151 U2 gnd 0.061857f
C152 P3 P1 0.009065f
C153 V2 m3_1120_n429# 1.87e-20
C154 MP P2 0.05668f
C155 G3 V3 0.055711f
C156 G2 V3 0.041965f
C157 NT G1 0.055711f
C158 C0 M0 0.055711f
C159 gnd AFF 0.127196f
C160 m2_1729_n327# L34 0.018008f
C161 vdd C4 0.094864f
C162 C3 vdd 0.094864f
C163 G2 m3_1120_n429# 0.004826f
C164 U3 L34 0.061857f
C165 OK OJ 0.058778f
C166 C2N U1 0.061857f
C167 vdd OJ 0.053537f
C168 A0 A0N1 1.62e-19
C169 gnd C4N 0.207735f
C170 V2 m2_1123_n465# 9.6e-20
C171 C2N m3_1054_n404# 1.12e-19
C172 P1 vdd 0.320929f
C173 Y0 B0 0.162736f
C174 C3N gnd 0.235227f
C175 HQ I2 0.05668f
C176 LO C1 0.055711f
C177 vdd P0 0.254168f
C178 G2 m2_1123_n465# 0.008947f
C179 U1 m2_937_n397# 9.6e-20
C180 KC KK 2.74e-19
C181 I0 vdd 0.149953f
C182 P1 P2 1.967832f
C183 KPK gnd 0.127196f
C184 B0N1 X0 4.82e-19
C185 C0 Z0 0.11336f
C186 vdd 6R 0.235619f
C187 C2 gnd 0.072183f
C188 C2N m2_937_n397# 0.018008f
C189 Y0 K0 0.055711f
C190 G2 m2_1729_n327# 6.24e-19
C191 P3 m3_1717_n374# 1.53e-19
C192 KP vdd 0.518157f
C193 U3 G2 0.041965f
C194 vdd X0 0.067556f
C195 P1 V1 0.056801f
C196 gnd AF 0.056518f
C197 KP P2 7.27e-19
C198 C1 UP 0.055711f
C199 GA gnd 0.092785f
C200 vdd m3_1054_n404# 0.001729f
C201 C4N C4 1.62e-19
C202 C3N C3 1.62e-19
C203 C2N vdd 0.06532f
C204 vdd m3_1717_n374# 0.003759f
C205 P3 vdd 0.365553f
C206 A0 m3_496_n300# 1.13e-19
C207 vdd m2_937_n397# 0.008839f
C208 I2 OJ 0.123714f
C209 B0N1 vdd 0.094864f
C210 I0 C3N 0.123714f
C211 V2 KC 0.247428f
C212 P3 P2 0.983916f
C213 U3 gnd 0.061857f
C214 vdd m2_453_n347# 0.00571f
C215 N0 gnd 0.061857f
C216 C2N V1 0.247428f
C217 C2N G1 0.055711f
C218 G2 KC 0.055711f
C219 OK vdd 0.194108f
C220 KPK I0 7.27e-19
C221 B0 N0 0.055711f
C222 A0 gnd 0.056518f
C223 G3 L34 0.055711f
C224 6R I2 7.27e-19
C225 G2 L34 0.174647f
C226 P1 AF 7.27e-19
C227 KP KPK 0.058778f
C228 GA P1 0.055711f
C229 m3_496_n300# A0N1 3.33e-19
C230 m2_937_n397# V1 9.6e-20
C231 KK gnd 0.127206f
C232 G1 m2_937_n397# 0.00987f
C233 A0 B0 0.227967f
C234 P1 m3_937_n361# 1.53e-19
C235 P2 vdd 0.449562f
C236 Z0 C1 0.11336f
C237 m2_496_n352# A0N1 2.88e-19
C238 C0 P0 0.241806f
C239 VE P1 0.05668f
C240 Z0 M0 0.061857f
C241 G2 V2 0.055711f
C242 gnd A0N1 0.072183f
C243 vdd V1 0.191129f
C244 U2 P2 0.041965f
C245 KK MP 3.8e-20
C246 G1 vdd 0.349941f
C247 KC gnd 0.118374f
C248 C2 m3_1054_n404# 1.87e-19
C249 HQ L34 2.74e-19
C250 OK AFF 0.135198f
C251 C2N C2 1.62e-19
C252 m3_1717_n374# V3 1.87e-20
C253 vdd AFF 0.147207f
C254 gnd L34 0.118374f
C255 m3_1503_n436# 0 0.01692f
C256 m3_1120_n429# 0 0.1404f
C257 m3_1054_n404# 0 0.016037f
C258 m3_2144_n302# 0 0.016037f
C259 m3_937_n361# 0 0.14305f
C260 m3_1717_n374# 0 0.120846f
C261 m3_496_n300# 0 0.084889f
C262 m2_1123_n465# 0 1.04973f
C263 m2_937_n397# 0 1.11581f
C264 m2_496_n352# 0 0.787321f
C265 m2_1729_n327# 0 0.666347f
C266 m2_453_n347# 0 1.7415f
C267 gnd 0 1.328833f **FLOATING
C268 N0 0 0.077618f **FLOATING
C269 vdd 0 43.72502f **FLOATING
C270 B0 0 1.061952f **FLOATING
C271 A0 0 1.339105f **FLOATING
C272 P2 0 1.980983f **FLOATING
C273 MP 0 0.080394f **FLOATING
C274 KK 0 0.869923f **FLOATING
C275 U2 0 0.079598f **FLOATING
C276 K0 0 0.077618f **FLOATING
C277 UP 0 0.054318f **FLOATING
C278 G1 0 1.318654f **FLOATING
C279 C3 0 0.019328f **FLOATING
C280 KC 0 0.556903f **FLOATING
C281 Y0 0 1.26094f **FLOATING
C282 P1 0 1.433693f **FLOATING
C283 C1 0 1.015367f **FLOATING
C284 C3N 0 0.380624f **FLOATING
C285 I0 0 0.067524f **FLOATING
C286 M0 0 0.077618f **FLOATING
C287 KPK 0 0.775747f **FLOATING
C288 KP 0 0.588774f **FLOATING
C289 V2 0 0.132907f **FLOATING
C290 C2 0 0.019328f **FLOATING
C291 U1 0 0.079598f **FLOATING
C292 G2 0 0.945851f **FLOATING
C293 GA 0 0.054318f **FLOATING
C294 C2N 0 0.556903f **FLOATING
C295 Z0 0 2.37156f **FLOATING
C296 C0 0 1.82639f **FLOATING
C297 P3 0 2.124685f **FLOATING
C298 AW 0 0.080394f **FLOATING
C299 VE 0 0.080394f **FLOATING
C300 B0N1 0 0.143763f **FLOATING
C301 HQ 0 0.83191f **FLOATING
C302 U3 0 0.079598f **FLOATING
C303 OK 0 0.939642f **FLOATING
C304 NT 0 0.054318f **FLOATING
C305 LO 0 0.054318f **FLOATING
C306 V1 0 0.132907f **FLOATING
C307 C4 0 0.019328f **FLOATING
C308 A0N1 0 0.041372f **FLOATING
C309 AFF 0 2.05566f **FLOATING
C310 OJ 0 0.383004f **FLOATING
C311 L34 0 0.556903f **FLOATING
C312 C4N 0 0.38067f **FLOATING
C313 P0 0 1.06873f **FLOATING
C314 I3 0 0.067524f **FLOATING
C315 I2 0 0.067524f **FLOATING
C316 6R 0 0.754516f **FLOATING
C317 LT 0 0.572436f **FLOATING
C318 V3 0 0.132907f **FLOATING
C319 X0 0 0.316742f **FLOATING
C320 G3 0 0.721943f **FLOATING
C321 AF 0 1.0581f **FLOATING
