magic
tech scmos
timestamp 1732052550
<< nwell >>
rect 742 -296 766 -278
rect 932 -289 956 -271
rect 831 -313 855 -295
rect 1021 -306 1045 -288
rect 1115 -292 1139 -274
rect 1318 -289 1342 -271
rect 1204 -309 1228 -291
rect 1407 -306 1431 -288
rect 742 -348 766 -330
rect 932 -341 956 -323
rect 1115 -344 1139 -326
rect 1318 -341 1342 -323
<< ntransistor >>
rect 812 -296 814 -290
rect 753 -307 755 -304
rect 1002 -289 1004 -283
rect 943 -300 945 -297
rect 1185 -292 1187 -286
rect 1126 -303 1128 -300
rect 1388 -289 1390 -283
rect 1329 -300 1331 -297
rect 1032 -317 1034 -314
rect 842 -324 844 -321
rect 1215 -320 1217 -317
rect 1418 -317 1420 -314
rect 812 -337 814 -331
rect 1002 -330 1004 -324
rect 1185 -333 1187 -327
rect 1388 -330 1390 -324
rect 943 -352 945 -349
rect 753 -359 755 -356
rect 1126 -355 1128 -352
rect 1329 -352 1331 -349
<< ptransistor >>
rect 943 -283 945 -277
rect 753 -290 755 -284
rect 1126 -286 1128 -280
rect 1329 -283 1331 -277
rect 1032 -300 1034 -294
rect 842 -307 844 -301
rect 1215 -303 1217 -297
rect 1418 -300 1420 -294
rect 753 -342 755 -336
rect 943 -335 945 -329
rect 1126 -338 1128 -332
rect 1329 -335 1331 -329
<< ndiffusion >>
rect 807 -296 812 -290
rect 814 -296 820 -290
rect 752 -307 753 -304
rect 755 -307 756 -304
rect 997 -289 1002 -283
rect 1004 -289 1010 -283
rect 942 -300 943 -297
rect 945 -300 946 -297
rect 1180 -292 1185 -286
rect 1187 -292 1193 -286
rect 1125 -303 1126 -300
rect 1128 -303 1129 -300
rect 1383 -289 1388 -283
rect 1390 -289 1396 -283
rect 1328 -300 1329 -297
rect 1331 -300 1332 -297
rect 1031 -317 1032 -314
rect 1034 -317 1035 -314
rect 841 -324 842 -321
rect 844 -324 845 -321
rect 1214 -320 1215 -317
rect 1217 -320 1218 -317
rect 1417 -317 1418 -314
rect 1420 -317 1421 -314
rect 808 -337 812 -331
rect 814 -337 820 -331
rect 998 -330 1002 -324
rect 1004 -330 1010 -324
rect 1181 -333 1185 -327
rect 1187 -333 1193 -327
rect 1384 -330 1388 -324
rect 1390 -330 1396 -324
rect 942 -352 943 -349
rect 945 -352 946 -349
rect 752 -359 753 -356
rect 755 -359 756 -356
rect 1125 -355 1126 -352
rect 1128 -355 1129 -352
rect 1328 -352 1329 -349
rect 1331 -352 1332 -349
<< pdiffusion >>
rect 942 -283 943 -277
rect 945 -283 946 -277
rect 752 -290 753 -284
rect 755 -290 756 -284
rect 1125 -286 1126 -280
rect 1128 -286 1129 -280
rect 1328 -283 1329 -277
rect 1331 -283 1332 -277
rect 1031 -300 1032 -294
rect 1034 -300 1035 -294
rect 841 -307 842 -301
rect 844 -307 845 -301
rect 1214 -303 1215 -297
rect 1217 -303 1218 -297
rect 1417 -300 1418 -294
rect 1420 -300 1421 -294
rect 752 -342 753 -336
rect 755 -342 756 -336
rect 942 -335 943 -329
rect 945 -335 946 -329
rect 1125 -338 1126 -332
rect 1128 -338 1129 -332
rect 1328 -335 1329 -329
rect 1331 -335 1332 -329
<< ndcontact >>
rect 803 -296 807 -290
rect 820 -296 824 -290
rect 748 -308 752 -304
rect 756 -307 760 -303
rect 993 -289 997 -283
rect 1010 -289 1014 -283
rect 938 -301 942 -297
rect 946 -300 950 -296
rect 1176 -292 1180 -286
rect 1193 -292 1197 -286
rect 1121 -304 1125 -300
rect 1129 -303 1133 -299
rect 1379 -289 1383 -283
rect 1396 -289 1400 -283
rect 1324 -301 1328 -297
rect 1332 -300 1336 -296
rect 1027 -318 1031 -314
rect 1035 -317 1039 -313
rect 837 -325 841 -321
rect 845 -324 849 -320
rect 1210 -321 1214 -317
rect 1218 -320 1222 -316
rect 1413 -318 1417 -314
rect 1421 -317 1425 -313
rect 803 -337 808 -331
rect 820 -337 824 -331
rect 993 -330 998 -324
rect 1010 -330 1014 -324
rect 1176 -333 1181 -327
rect 1193 -333 1197 -327
rect 1379 -330 1384 -324
rect 1396 -330 1400 -324
rect 938 -353 942 -349
rect 946 -352 950 -348
rect 748 -360 752 -356
rect 756 -359 760 -355
rect 1121 -356 1125 -352
rect 1129 -355 1133 -351
rect 1324 -353 1328 -349
rect 1332 -352 1336 -348
<< pdcontact >>
rect 938 -283 942 -277
rect 946 -283 950 -277
rect 748 -290 752 -284
rect 756 -290 760 -284
rect 1121 -286 1125 -280
rect 1129 -286 1133 -280
rect 1324 -283 1328 -277
rect 1332 -283 1336 -277
rect 1027 -300 1031 -294
rect 1035 -300 1039 -294
rect 837 -307 841 -301
rect 845 -307 849 -301
rect 1210 -303 1214 -297
rect 1218 -303 1222 -297
rect 1413 -300 1417 -294
rect 1421 -300 1425 -294
rect 748 -342 752 -336
rect 756 -342 760 -336
rect 938 -335 942 -329
rect 946 -335 950 -329
rect 1121 -338 1125 -332
rect 1129 -338 1133 -332
rect 1324 -335 1328 -329
rect 1332 -335 1336 -329
<< polysilicon >>
rect 943 -277 945 -274
rect 1329 -277 1331 -274
rect 753 -284 755 -281
rect 1126 -280 1128 -277
rect 1002 -283 1004 -280
rect 812 -290 814 -287
rect 753 -304 755 -290
rect 812 -305 814 -296
rect 943 -297 945 -283
rect 1388 -283 1390 -280
rect 1185 -286 1187 -283
rect 842 -301 844 -298
rect 1002 -298 1004 -289
rect 1032 -294 1034 -291
rect 1126 -300 1128 -286
rect 943 -303 945 -300
rect 753 -310 755 -307
rect 842 -321 844 -307
rect 1032 -314 1034 -300
rect 1185 -301 1187 -292
rect 1215 -297 1217 -294
rect 1329 -297 1331 -283
rect 1388 -298 1390 -289
rect 1418 -294 1420 -291
rect 1329 -303 1331 -300
rect 1126 -306 1128 -303
rect 1215 -317 1217 -303
rect 1418 -314 1420 -300
rect 1032 -320 1034 -317
rect 1418 -320 1420 -317
rect 1002 -324 1004 -321
rect 1215 -323 1217 -320
rect 1388 -324 1390 -321
rect 842 -327 844 -324
rect 812 -331 814 -328
rect 943 -329 945 -326
rect 753 -336 755 -333
rect 1185 -327 1187 -324
rect 753 -349 755 -342
rect 812 -346 814 -337
rect 943 -342 945 -335
rect 1002 -339 1004 -330
rect 1126 -332 1128 -329
rect 1329 -329 1331 -326
rect 942 -346 945 -342
rect 1126 -345 1128 -338
rect 1185 -342 1187 -333
rect 1329 -342 1331 -335
rect 1388 -339 1390 -330
rect 943 -349 945 -346
rect 752 -353 755 -349
rect 1125 -349 1128 -345
rect 1328 -346 1331 -342
rect 1329 -349 1331 -346
rect 1126 -352 1128 -349
rect 753 -356 755 -353
rect 943 -355 945 -352
rect 1329 -355 1331 -352
rect 1126 -358 1128 -355
rect 753 -362 755 -359
<< polycontact >>
rect 749 -301 753 -297
rect 939 -294 943 -290
rect 808 -305 812 -300
rect 998 -298 1002 -293
rect 1122 -297 1126 -293
rect 838 -318 842 -314
rect 1028 -311 1032 -307
rect 1181 -301 1185 -296
rect 1325 -294 1329 -290
rect 1384 -298 1388 -293
rect 1211 -314 1215 -310
rect 1414 -311 1418 -307
rect 808 -346 812 -342
rect 998 -339 1002 -335
rect 938 -346 942 -342
rect 1181 -342 1185 -338
rect 1384 -339 1388 -335
rect 748 -353 752 -349
rect 1121 -349 1125 -345
rect 1324 -346 1328 -342
<< metal1 >>
rect 923 -263 997 -258
rect 733 -270 807 -265
rect 733 -297 737 -270
rect 742 -279 766 -275
rect 748 -284 752 -279
rect 803 -290 807 -270
rect 923 -290 927 -263
rect 932 -272 956 -268
rect 938 -277 942 -272
rect 993 -283 997 -263
rect 1106 -266 1180 -261
rect 1021 -289 1045 -285
rect 831 -296 855 -292
rect 908 -294 939 -290
rect 723 -301 749 -297
rect 748 -311 752 -308
rect 742 -315 766 -311
rect 820 -314 824 -296
rect 837 -301 841 -296
rect 938 -304 942 -301
rect 932 -308 956 -304
rect 1010 -307 1014 -289
rect 1027 -294 1031 -289
rect 1106 -293 1110 -266
rect 1115 -275 1139 -271
rect 1121 -280 1125 -275
rect 1176 -286 1180 -266
rect 1309 -263 1383 -258
rect 1204 -292 1228 -288
rect 1309 -290 1313 -263
rect 1318 -272 1342 -268
rect 1324 -277 1328 -272
rect 1379 -283 1383 -263
rect 1407 -289 1431 -285
rect 1095 -297 1122 -293
rect 1121 -307 1125 -304
rect 1010 -311 1028 -307
rect 1115 -311 1139 -307
rect 1193 -310 1197 -292
rect 1210 -297 1214 -292
rect 1300 -294 1325 -290
rect 1324 -304 1328 -301
rect 1318 -308 1342 -304
rect 1396 -307 1400 -289
rect 1413 -294 1417 -289
rect 820 -318 838 -314
rect 742 -331 766 -327
rect 820 -331 824 -318
rect 932 -324 956 -320
rect 1010 -324 1014 -311
rect 1193 -314 1211 -310
rect 1396 -311 1414 -307
rect 1027 -321 1031 -318
rect 837 -328 841 -325
rect 748 -336 752 -331
rect 831 -332 855 -328
rect 938 -329 942 -324
rect 1021 -325 1045 -321
rect 1115 -327 1139 -323
rect 1193 -327 1197 -314
rect 1210 -324 1214 -321
rect 1318 -324 1342 -320
rect 1396 -324 1400 -311
rect 1413 -321 1417 -318
rect 1121 -332 1125 -327
rect 1204 -328 1228 -324
rect 1324 -329 1328 -324
rect 1407 -325 1431 -321
rect 938 -356 942 -353
rect 1324 -356 1328 -353
rect 932 -360 956 -356
rect 1121 -359 1125 -356
rect 748 -363 752 -360
rect 1115 -363 1139 -359
rect 1318 -360 1342 -356
rect 742 -367 766 -363
<< metal2 >>
rect 986 -298 998 -293
rect 796 -305 808 -300
rect 796 -320 800 -305
rect 986 -313 990 -298
rect 734 -324 800 -320
rect 924 -317 990 -313
rect 1169 -301 1181 -296
rect 1372 -298 1384 -293
rect 1169 -316 1173 -301
rect 1372 -313 1376 -298
rect 734 -346 738 -324
rect 924 -339 928 -317
rect 1107 -320 1173 -316
rect 1310 -317 1376 -313
rect 908 -342 928 -339
rect 946 -342 950 -335
rect 989 -339 998 -335
rect 989 -342 993 -339
rect 1107 -342 1111 -320
rect 723 -349 738 -346
rect 756 -349 760 -342
rect 799 -346 808 -342
rect 908 -343 938 -342
rect 924 -346 938 -343
rect 946 -346 993 -342
rect 1095 -345 1111 -342
rect 1129 -345 1133 -338
rect 1172 -342 1181 -338
rect 1310 -339 1314 -317
rect 1300 -342 1314 -339
rect 1332 -342 1336 -335
rect 1375 -339 1384 -335
rect 1375 -342 1379 -339
rect 1172 -345 1176 -342
rect 1300 -343 1324 -342
rect 1095 -346 1121 -345
rect 799 -349 803 -346
rect 946 -348 950 -346
rect 1107 -349 1121 -346
rect 1129 -349 1176 -345
rect 1310 -346 1324 -343
rect 1332 -346 1379 -342
rect 1332 -348 1336 -346
rect 723 -350 748 -349
rect 734 -353 748 -350
rect 756 -353 803 -349
rect 1129 -351 1133 -349
rect 756 -355 760 -353
<< metal3 >>
rect 946 -289 950 -283
rect 756 -296 760 -290
rect 946 -294 978 -289
rect 946 -296 950 -294
rect 756 -301 788 -296
rect 756 -303 760 -301
rect 784 -331 788 -301
rect 845 -314 849 -307
rect 845 -318 855 -314
rect 845 -320 849 -318
rect 974 -324 978 -294
rect 1129 -292 1133 -286
rect 1332 -289 1336 -283
rect 1129 -297 1161 -292
rect 1332 -294 1364 -289
rect 1332 -296 1336 -294
rect 1129 -299 1133 -297
rect 1035 -307 1039 -300
rect 1035 -311 1045 -307
rect 1035 -313 1039 -311
rect 974 -330 993 -324
rect 1157 -327 1161 -297
rect 1218 -310 1222 -303
rect 1218 -314 1228 -310
rect 1218 -316 1222 -314
rect 1360 -324 1364 -294
rect 1421 -307 1425 -300
rect 1421 -311 1431 -307
rect 1421 -313 1425 -311
rect 784 -337 803 -331
rect 1157 -333 1176 -327
rect 1360 -330 1379 -324
<< labels >>
rlabel nwell 762 -282 764 -280 1 vdd
rlabel pdcontact 748 -290 752 -284 1 vdd
rlabel nwell 762 -334 764 -332 1 vdd
rlabel pdcontact 748 -342 752 -336 1 vdd
rlabel nwell 851 -299 853 -297 1 vdd
rlabel pdcontact 837 -307 841 -301 1 vdd
rlabel ndcontact 837 -325 841 -321 1 gnd
rlabel ndcontact 748 -308 752 -304 1 gnd
rlabel ndcontact 748 -360 752 -356 1 gnd
rlabel polycontact 749 -301 753 -297 1 P0
rlabel polycontact 748 -353 752 -349 1 C0
rlabel polycontact 808 -305 812 -300 1 C0
rlabel ndcontact 756 -307 760 -303 1 P0N1
rlabel ndcontact 803 -337 807 -332 1 P0N1
rlabel pdcontact 756 -342 760 -336 1 C0N1
rlabel ndcontact 756 -359 760 -355 1 C0N1
rlabel polycontact 808 -346 812 -342 1 C0N1
rlabel ndcontact 803 -296 807 -291 1 P0
rlabel ndcontact 820 -295 824 -291 1 S0N
rlabel ndcontact 820 -336 824 -332 1 S0N
rlabel polycontact 838 -318 842 -314 1 S0N
rlabel ndcontact 845 -324 849 -320 1 S0
rlabel pdcontact 845 -307 849 -301 1 S0
rlabel pdcontact 756 -290 760 -284 1 P0N1
rlabel nwell 952 -275 954 -273 1 vdd
rlabel pdcontact 938 -283 942 -277 1 vdd
rlabel nwell 952 -327 954 -325 1 vdd
rlabel pdcontact 938 -335 942 -329 1 vdd
rlabel nwell 1041 -292 1043 -290 1 vdd
rlabel pdcontact 1027 -300 1031 -294 1 vdd
rlabel ndcontact 1027 -318 1031 -314 1 gnd
rlabel ndcontact 938 -301 942 -297 1 gnd
rlabel ndcontact 938 -353 942 -349 1 gnd
rlabel polycontact 939 -294 943 -290 1 P1
rlabel polycontact 938 -346 942 -342 1 C1
rlabel pdcontact 946 -335 950 -329 1 C1N1
rlabel ndcontact 946 -352 950 -348 1 C1N1
rlabel polycontact 998 -339 1002 -335 1 C1N1
rlabel ndcontact 946 -300 950 -296 1 P1N1
rlabel pdcontact 946 -283 950 -277 1 P1N1
rlabel ndcontact 993 -330 997 -325 1 P1N1
rlabel polycontact 998 -298 1002 -293 1 C1
rlabel ndcontact 1010 -329 1014 -325 1 S1N
rlabel ndcontact 1010 -288 1014 -284 1 S1N
rlabel polycontact 1028 -311 1032 -307 1 S1N
rlabel ndcontact 1035 -317 1039 -313 1 S1
rlabel pdcontact 1035 -300 1039 -294 1 S1
rlabel ndcontact 993 -289 997 -283 1 P1
rlabel nwell 1135 -278 1137 -276 1 vdd
rlabel pdcontact 1121 -286 1125 -280 1 vdd
rlabel nwell 1135 -330 1137 -328 1 vdd
rlabel pdcontact 1121 -338 1125 -332 1 vdd
rlabel nwell 1224 -295 1226 -293 1 vdd
rlabel pdcontact 1210 -303 1214 -297 1 vdd
rlabel ndcontact 1210 -321 1214 -317 1 gnd
rlabel ndcontact 1121 -304 1125 -300 1 gnd
rlabel ndcontact 1121 -356 1125 -352 1 gnd
rlabel polycontact 1122 -297 1126 -293 1 P2
rlabel ndcontact 1129 -303 1133 -299 1 P2N1
rlabel pdcontact 1129 -286 1133 -280 1 P2N1
rlabel ndcontact 1176 -333 1180 -327 1 P2N1
rlabel polycontact 1121 -349 1125 -345 1 C2
rlabel pdcontact 1129 -338 1133 -332 1 C2N1
rlabel ndcontact 1129 -355 1133 -351 1 C2N1
rlabel polycontact 1181 -342 1185 -338 1 C2N1
rlabel polycontact 1181 -301 1185 -296 1 C2
rlabel ndcontact 1193 -332 1197 -327 1 S2N
rlabel ndcontact 1193 -291 1197 -286 1 S2N
rlabel polycontact 1211 -314 1215 -310 1 S2N
rlabel pdcontact 1218 -303 1222 -297 1 S2
rlabel ndcontact 1218 -320 1222 -316 1 S2
rlabel nwell 1338 -275 1340 -273 1 vdd
rlabel pdcontact 1324 -283 1328 -277 1 vdd
rlabel nwell 1338 -327 1340 -325 1 vdd
rlabel pdcontact 1324 -335 1328 -329 1 vdd
rlabel nwell 1427 -292 1429 -290 1 vdd
rlabel pdcontact 1413 -300 1417 -294 1 vdd
rlabel ndcontact 1413 -318 1417 -314 1 gnd
rlabel ndcontact 1324 -301 1328 -297 1 gnd
rlabel ndcontact 1324 -353 1328 -349 1 gnd
rlabel polycontact 1325 -294 1329 -290 1 P3
rlabel ndcontact 1332 -300 1336 -296 1 P3N1
rlabel pdcontact 1332 -283 1336 -277 1 P3N1
rlabel ndcontact 1379 -330 1383 -324 1 P3N1
rlabel polycontact 1324 -346 1328 -342 1 C3
rlabel pdcontact 1332 -335 1336 -329 1 C3N1
rlabel ndcontact 1332 -352 1336 -348 1 C3N1
rlabel polycontact 1384 -339 1388 -335 1 C3N1
rlabel polycontact 1384 -298 1388 -293 1 C3
rlabel ndcontact 1379 -289 1383 -283 1 P3
rlabel ndcontact 1396 -329 1400 -324 1 S3N
rlabel ndcontact 1396 -288 1400 -283 1 S3N
rlabel polycontact 1414 -311 1418 -307 1 S3N
rlabel ndcontact 1421 -317 1425 -313 1 S3
rlabel pdcontact 1421 -300 1425 -294 1 S3
rlabel ndcontact 1176 -292 1180 -286 1 P2
<< end >>
