magic
tech scmos
timestamp 1732051050
<< nwell >>
rect 1409 -247 1433 -229
rect 1498 -264 1522 -246
rect 1669 -250 1693 -232
rect 1758 -267 1782 -249
rect 482 -293 506 -275
rect 571 -310 595 -292
rect 651 -296 675 -278
rect 716 -313 740 -295
rect 1409 -299 1433 -281
rect 1669 -302 1693 -284
rect 482 -345 506 -327
rect 651 -348 675 -330
rect 988 -357 1012 -339
rect 587 -396 647 -362
rect 1063 -374 1087 -356
rect 1133 -360 1157 -342
rect 1222 -377 1246 -359
rect 1404 -369 1464 -335
rect 988 -409 1012 -391
rect 1133 -412 1157 -394
rect 1459 -401 1483 -383
rect 665 -453 725 -419
rect 1568 -422 1654 -340
rect 1686 -427 1747 -365
rect 1809 -414 1878 -354
rect 1887 -414 1911 -396
rect 983 -479 1043 -445
rect 588 -532 648 -498
rect 1038 -511 1062 -493
rect 1103 -499 1164 -437
rect 1753 -440 1777 -422
rect 1940 -423 1965 -366
rect 1986 -411 2010 -393
rect 2052 -423 2077 -366
rect 2092 -408 2116 -390
rect 1170 -512 1194 -494
rect 1647 -526 1671 -508
rect 1040 -706 1064 -688
rect 1129 -723 1153 -705
rect 1300 -709 1324 -691
rect 1389 -726 1413 -708
rect 1040 -758 1064 -740
rect 1300 -761 1324 -743
rect 1035 -822 1095 -788
rect 1090 -854 1114 -836
rect 1179 -861 1240 -799
rect 1336 -848 1405 -788
rect 1246 -874 1270 -856
rect 1445 -857 1470 -800
<< ntransistor >>
rect 1479 -247 1481 -241
rect 1420 -258 1422 -255
rect 1739 -250 1741 -244
rect 1680 -261 1682 -258
rect 1509 -275 1511 -272
rect 1769 -278 1771 -275
rect 552 -293 554 -287
rect 493 -304 495 -301
rect 697 -296 699 -290
rect 1479 -288 1481 -282
rect 662 -307 664 -304
rect 1739 -291 1741 -285
rect 582 -321 584 -318
rect 1420 -310 1422 -307
rect 1680 -313 1682 -310
rect 727 -324 729 -321
rect 552 -334 554 -328
rect 697 -337 699 -331
rect 493 -356 495 -353
rect 662 -359 664 -356
rect 1044 -357 1046 -351
rect 999 -368 1001 -365
rect 1203 -360 1205 -354
rect 1144 -371 1146 -368
rect 1074 -385 1076 -382
rect 1233 -388 1235 -385
rect 1044 -398 1046 -392
rect 1203 -401 1205 -395
rect 1433 -396 1435 -390
rect 1470 -412 1472 -409
rect 616 -423 618 -417
rect 999 -420 1001 -417
rect 1144 -423 1146 -420
rect 1433 -422 1435 -416
rect 1898 -425 1900 -422
rect 1997 -422 1999 -419
rect 2103 -419 2105 -416
rect 616 -449 618 -443
rect 1607 -447 1609 -438
rect 1848 -439 1850 -430
rect 1962 -440 1964 -434
rect 1944 -447 1946 -441
rect 2074 -440 2076 -434
rect 2056 -447 2058 -441
rect 1727 -454 1729 -448
rect 1764 -451 1766 -448
rect 1607 -467 1609 -458
rect 1848 -459 1850 -450
rect 1704 -467 1706 -461
rect 694 -480 696 -474
rect 1727 -480 1729 -474
rect 1607 -495 1609 -486
rect 1848 -487 1850 -478
rect 694 -506 696 -500
rect 1012 -506 1014 -500
rect 1049 -522 1051 -519
rect 1607 -515 1609 -506
rect 1144 -526 1146 -520
rect 1181 -523 1183 -520
rect 1012 -532 1014 -526
rect 1121 -539 1123 -533
rect 1658 -537 1660 -534
rect 1144 -552 1146 -546
rect 617 -559 619 -553
rect 617 -585 619 -579
rect 1110 -706 1112 -700
rect 1051 -717 1053 -714
rect 1370 -709 1372 -703
rect 1311 -720 1313 -717
rect 1140 -734 1142 -731
rect 1400 -737 1402 -734
rect 1110 -747 1112 -741
rect 1370 -750 1372 -744
rect 1051 -769 1053 -766
rect 1311 -772 1313 -769
rect 1064 -849 1066 -843
rect 1101 -865 1103 -862
rect 1064 -875 1066 -869
rect 1375 -873 1377 -864
rect 1467 -874 1469 -868
rect 1449 -881 1451 -875
rect 1220 -888 1222 -882
rect 1257 -885 1259 -882
rect 1375 -893 1377 -884
rect 1197 -901 1199 -895
rect 1220 -914 1222 -908
rect 1375 -921 1377 -912
<< ptransistor >>
rect 1420 -241 1422 -235
rect 1680 -244 1682 -238
rect 1509 -258 1511 -252
rect 1769 -261 1771 -255
rect 493 -287 495 -281
rect 662 -290 664 -284
rect 582 -304 584 -298
rect 1420 -293 1422 -287
rect 1680 -296 1682 -290
rect 727 -307 729 -301
rect 493 -339 495 -333
rect 662 -342 664 -336
rect 999 -351 1001 -345
rect 1425 -347 1427 -341
rect 1144 -354 1146 -348
rect 608 -374 610 -368
rect 1074 -368 1076 -362
rect 1451 -363 1453 -357
rect 1640 -361 1642 -349
rect 1233 -371 1235 -365
rect 634 -390 636 -384
rect 1623 -381 1625 -369
rect 999 -403 1001 -397
rect 1144 -406 1146 -400
rect 1470 -395 1472 -389
rect 1603 -395 1605 -383
rect 1711 -385 1713 -373
rect 1864 -373 1866 -361
rect 1844 -387 1846 -375
rect 1952 -384 1954 -372
rect 2064 -384 2066 -372
rect 1584 -413 1586 -401
rect 1825 -405 1827 -393
rect 1703 -419 1705 -407
rect 1734 -419 1736 -407
rect 1898 -408 1900 -402
rect 686 -431 688 -425
rect 1952 -416 1954 -404
rect 1997 -405 1999 -399
rect 2103 -402 2105 -396
rect 2064 -416 2066 -404
rect 1764 -434 1766 -428
rect 712 -447 714 -441
rect 1004 -457 1006 -451
rect 1128 -457 1130 -445
rect 1030 -473 1032 -467
rect 1120 -491 1122 -479
rect 1151 -491 1153 -479
rect 609 -510 611 -504
rect 1049 -505 1051 -499
rect 1181 -506 1183 -500
rect 635 -526 637 -520
rect 1658 -520 1660 -514
rect 1051 -700 1053 -694
rect 1311 -703 1313 -697
rect 1140 -717 1142 -711
rect 1400 -720 1402 -714
rect 1051 -752 1053 -746
rect 1311 -755 1313 -749
rect 1056 -800 1058 -794
rect 1082 -816 1084 -810
rect 1204 -819 1206 -807
rect 1391 -807 1393 -795
rect 1371 -821 1373 -809
rect 1457 -818 1459 -806
rect 1352 -839 1354 -827
rect 1101 -848 1103 -842
rect 1196 -853 1198 -841
rect 1227 -853 1229 -841
rect 1457 -850 1459 -838
rect 1257 -868 1259 -862
<< ndiffusion >>
rect 1474 -247 1479 -241
rect 1481 -247 1487 -241
rect 1419 -258 1420 -255
rect 1422 -258 1423 -255
rect 1734 -250 1739 -244
rect 1741 -250 1747 -244
rect 1679 -261 1680 -258
rect 1682 -261 1683 -258
rect 1508 -275 1509 -272
rect 1511 -275 1512 -272
rect 1768 -278 1769 -275
rect 1771 -278 1772 -275
rect 547 -293 552 -287
rect 554 -293 560 -287
rect 492 -304 493 -301
rect 495 -304 496 -301
rect 692 -296 697 -290
rect 699 -296 705 -290
rect 1475 -288 1479 -282
rect 1481 -288 1487 -282
rect 661 -307 662 -304
rect 664 -307 665 -304
rect 1735 -291 1739 -285
rect 1741 -291 1747 -285
rect 581 -321 582 -318
rect 584 -321 585 -318
rect 1419 -310 1420 -307
rect 1422 -310 1423 -307
rect 1679 -313 1680 -310
rect 1682 -313 1683 -310
rect 726 -324 727 -321
rect 729 -324 730 -321
rect 548 -334 552 -328
rect 554 -334 560 -328
rect 693 -337 697 -331
rect 699 -337 705 -331
rect 492 -356 493 -353
rect 495 -356 496 -353
rect 661 -359 662 -356
rect 664 -359 665 -356
rect 1039 -357 1044 -351
rect 1046 -357 1052 -351
rect 998 -368 999 -365
rect 1001 -368 1002 -365
rect 1198 -360 1203 -354
rect 1205 -360 1211 -354
rect 1143 -371 1144 -368
rect 1146 -371 1147 -368
rect 1073 -385 1074 -382
rect 1076 -385 1077 -382
rect 1232 -388 1233 -385
rect 1235 -388 1236 -385
rect 1040 -398 1044 -392
rect 1046 -398 1052 -392
rect 1199 -401 1203 -395
rect 1205 -401 1211 -395
rect 1432 -396 1433 -390
rect 1435 -396 1436 -390
rect 1469 -412 1470 -409
rect 1472 -412 1473 -409
rect 615 -423 616 -417
rect 618 -423 619 -417
rect 998 -420 999 -417
rect 1001 -420 1002 -417
rect 1143 -423 1144 -420
rect 1146 -423 1147 -420
rect 1432 -422 1433 -416
rect 1435 -422 1436 -416
rect 1897 -425 1898 -422
rect 1900 -425 1901 -422
rect 1996 -422 1997 -419
rect 1999 -422 2000 -419
rect 2102 -419 2103 -416
rect 2105 -419 2106 -416
rect 615 -449 616 -443
rect 618 -449 619 -443
rect 1606 -447 1607 -438
rect 1609 -447 1610 -438
rect 1847 -439 1848 -430
rect 1850 -439 1851 -430
rect 1961 -440 1962 -434
rect 1964 -440 1965 -434
rect 1943 -447 1944 -441
rect 1946 -447 1947 -441
rect 2073 -440 2074 -434
rect 2076 -440 2077 -434
rect 2055 -447 2056 -441
rect 2058 -447 2059 -441
rect 1726 -454 1727 -448
rect 1729 -454 1730 -448
rect 1763 -451 1764 -448
rect 1766 -451 1767 -448
rect 1606 -467 1607 -458
rect 1609 -467 1610 -458
rect 1847 -459 1848 -450
rect 1850 -459 1851 -450
rect 1703 -467 1704 -461
rect 1706 -467 1707 -461
rect 693 -480 694 -474
rect 696 -480 697 -474
rect 1726 -480 1727 -474
rect 1729 -480 1730 -474
rect 1606 -495 1607 -486
rect 1609 -495 1610 -486
rect 1847 -487 1848 -478
rect 1850 -487 1851 -478
rect 693 -506 694 -500
rect 696 -506 697 -500
rect 1011 -506 1012 -500
rect 1014 -506 1015 -500
rect 1048 -522 1049 -519
rect 1051 -522 1052 -519
rect 1606 -515 1607 -506
rect 1609 -515 1610 -506
rect 1143 -526 1144 -520
rect 1146 -526 1147 -520
rect 1180 -523 1181 -520
rect 1183 -523 1184 -520
rect 1011 -532 1012 -526
rect 1014 -532 1015 -526
rect 1120 -539 1121 -533
rect 1123 -539 1124 -533
rect 1657 -537 1658 -534
rect 1660 -537 1661 -534
rect 1143 -552 1144 -546
rect 1146 -552 1147 -546
rect 616 -559 617 -553
rect 619 -559 620 -553
rect 616 -585 617 -579
rect 619 -585 620 -579
rect 1105 -706 1110 -700
rect 1112 -706 1118 -700
rect 1050 -717 1051 -714
rect 1053 -717 1054 -714
rect 1365 -709 1370 -703
rect 1372 -709 1378 -703
rect 1310 -720 1311 -717
rect 1313 -720 1314 -717
rect 1139 -734 1140 -731
rect 1142 -734 1143 -731
rect 1399 -737 1400 -734
rect 1402 -737 1403 -734
rect 1106 -747 1110 -741
rect 1112 -747 1118 -741
rect 1366 -750 1370 -744
rect 1372 -750 1378 -744
rect 1050 -769 1051 -766
rect 1053 -769 1054 -766
rect 1310 -772 1311 -769
rect 1313 -772 1314 -769
rect 1063 -849 1064 -843
rect 1066 -849 1067 -843
rect 1100 -865 1101 -862
rect 1103 -865 1104 -862
rect 1063 -875 1064 -869
rect 1066 -875 1067 -869
rect 1374 -873 1375 -864
rect 1377 -873 1378 -864
rect 1466 -874 1467 -868
rect 1469 -874 1470 -868
rect 1448 -881 1449 -875
rect 1451 -881 1452 -875
rect 1219 -888 1220 -882
rect 1222 -888 1223 -882
rect 1256 -885 1257 -882
rect 1259 -885 1260 -882
rect 1374 -893 1375 -884
rect 1377 -893 1378 -884
rect 1196 -901 1197 -895
rect 1199 -901 1200 -895
rect 1219 -914 1220 -908
rect 1222 -914 1223 -908
rect 1374 -921 1375 -912
rect 1377 -921 1378 -912
<< pdiffusion >>
rect 1419 -241 1420 -235
rect 1422 -241 1423 -235
rect 1679 -244 1680 -238
rect 1682 -244 1683 -238
rect 1508 -258 1509 -252
rect 1511 -258 1512 -252
rect 1768 -261 1769 -255
rect 1771 -261 1772 -255
rect 492 -287 493 -281
rect 495 -287 496 -281
rect 661 -290 662 -284
rect 664 -290 665 -284
rect 581 -304 582 -298
rect 584 -304 585 -298
rect 1419 -293 1420 -287
rect 1422 -293 1423 -287
rect 1679 -296 1680 -290
rect 1682 -296 1683 -290
rect 726 -307 727 -301
rect 729 -307 730 -301
rect 492 -339 493 -333
rect 495 -339 496 -333
rect 661 -342 662 -336
rect 664 -342 665 -336
rect 998 -351 999 -345
rect 1001 -351 1002 -345
rect 1424 -347 1425 -341
rect 1427 -347 1428 -341
rect 1143 -354 1144 -348
rect 1146 -354 1147 -348
rect 607 -374 608 -368
rect 610 -374 611 -368
rect 1073 -368 1074 -362
rect 1076 -368 1077 -362
rect 1450 -363 1451 -357
rect 1453 -363 1454 -357
rect 1639 -361 1640 -349
rect 1642 -361 1643 -349
rect 1232 -371 1233 -365
rect 1235 -371 1236 -365
rect 633 -390 634 -384
rect 636 -390 637 -384
rect 1622 -381 1623 -369
rect 1625 -381 1626 -369
rect 998 -403 999 -397
rect 1001 -403 1002 -397
rect 1143 -406 1144 -400
rect 1146 -406 1147 -400
rect 1469 -395 1470 -389
rect 1472 -395 1473 -389
rect 1602 -395 1603 -383
rect 1605 -395 1606 -383
rect 1710 -385 1711 -373
rect 1713 -385 1714 -373
rect 1863 -373 1864 -361
rect 1866 -373 1867 -361
rect 1843 -387 1844 -375
rect 1846 -387 1847 -375
rect 1951 -384 1952 -372
rect 1954 -384 1955 -372
rect 2063 -384 2064 -372
rect 2066 -384 2067 -372
rect 1583 -413 1584 -401
rect 1586 -413 1587 -401
rect 1824 -405 1825 -393
rect 1827 -405 1828 -393
rect 1702 -419 1703 -407
rect 1705 -419 1706 -407
rect 1733 -419 1734 -407
rect 1736 -419 1737 -407
rect 1897 -408 1898 -402
rect 1900 -408 1901 -402
rect 685 -431 686 -425
rect 688 -431 689 -425
rect 1951 -416 1952 -404
rect 1954 -416 1955 -404
rect 1996 -405 1997 -399
rect 1999 -405 2000 -399
rect 2102 -402 2103 -396
rect 2105 -402 2106 -396
rect 2063 -416 2064 -404
rect 2066 -416 2067 -404
rect 1763 -434 1764 -428
rect 1766 -434 1767 -428
rect 711 -447 712 -441
rect 714 -447 715 -441
rect 1003 -457 1004 -451
rect 1006 -457 1007 -451
rect 1127 -457 1128 -445
rect 1130 -457 1131 -445
rect 1029 -473 1030 -467
rect 1032 -473 1033 -467
rect 1119 -491 1120 -479
rect 1122 -491 1123 -479
rect 1150 -491 1151 -479
rect 1153 -491 1154 -479
rect 608 -510 609 -504
rect 611 -510 612 -504
rect 1048 -505 1049 -499
rect 1051 -505 1052 -499
rect 1180 -506 1181 -500
rect 1183 -506 1184 -500
rect 634 -526 635 -520
rect 637 -526 638 -520
rect 1657 -520 1658 -514
rect 1660 -520 1661 -514
rect 1050 -700 1051 -694
rect 1053 -700 1054 -694
rect 1310 -703 1311 -697
rect 1313 -703 1314 -697
rect 1139 -717 1140 -711
rect 1142 -717 1143 -711
rect 1399 -720 1400 -714
rect 1402 -720 1403 -714
rect 1050 -752 1051 -746
rect 1053 -752 1054 -746
rect 1310 -755 1311 -749
rect 1313 -755 1314 -749
rect 1055 -800 1056 -794
rect 1058 -800 1059 -794
rect 1081 -816 1082 -810
rect 1084 -816 1085 -810
rect 1203 -819 1204 -807
rect 1206 -819 1207 -807
rect 1390 -807 1391 -795
rect 1393 -807 1394 -795
rect 1370 -821 1371 -809
rect 1373 -821 1374 -809
rect 1456 -818 1457 -806
rect 1459 -818 1460 -806
rect 1351 -839 1352 -827
rect 1354 -839 1355 -827
rect 1100 -848 1101 -842
rect 1103 -848 1104 -842
rect 1195 -853 1196 -841
rect 1198 -853 1199 -841
rect 1226 -853 1227 -841
rect 1229 -853 1230 -841
rect 1456 -850 1457 -838
rect 1459 -850 1460 -838
rect 1256 -868 1257 -862
rect 1259 -868 1260 -862
<< ndcontact >>
rect 1470 -247 1474 -241
rect 1487 -247 1491 -241
rect 1415 -259 1419 -255
rect 1423 -258 1427 -254
rect 1730 -250 1734 -244
rect 1747 -250 1751 -244
rect 1675 -262 1679 -258
rect 1683 -261 1687 -257
rect 1504 -276 1508 -272
rect 1512 -275 1516 -271
rect 1764 -279 1768 -275
rect 1772 -278 1776 -274
rect 543 -293 547 -287
rect 560 -293 564 -287
rect 488 -305 492 -301
rect 496 -304 500 -300
rect 688 -296 692 -290
rect 705 -296 709 -290
rect 1470 -288 1475 -282
rect 1487 -288 1491 -282
rect 657 -308 661 -304
rect 665 -307 669 -303
rect 1730 -291 1735 -285
rect 1747 -291 1751 -285
rect 577 -322 581 -318
rect 585 -321 589 -317
rect 1415 -311 1419 -307
rect 1423 -310 1427 -306
rect 1675 -314 1679 -310
rect 1683 -313 1687 -309
rect 722 -325 726 -321
rect 730 -324 734 -320
rect 543 -334 548 -328
rect 560 -334 564 -328
rect 688 -337 693 -331
rect 705 -337 709 -331
rect 488 -357 492 -353
rect 496 -356 500 -352
rect 657 -360 661 -356
rect 665 -359 669 -355
rect 1035 -357 1039 -351
rect 1052 -357 1056 -351
rect 994 -369 998 -365
rect 1002 -368 1006 -364
rect 1194 -360 1198 -354
rect 1211 -360 1215 -354
rect 1139 -372 1143 -368
rect 1147 -371 1151 -367
rect 1069 -386 1073 -382
rect 1077 -385 1081 -381
rect 1228 -389 1232 -385
rect 1236 -388 1240 -384
rect 1035 -398 1040 -392
rect 1052 -398 1056 -392
rect 1194 -401 1199 -395
rect 1211 -401 1215 -395
rect 1428 -396 1432 -390
rect 1436 -396 1440 -390
rect 1465 -413 1469 -409
rect 1473 -412 1477 -408
rect 611 -423 615 -417
rect 619 -423 623 -417
rect 994 -421 998 -417
rect 1002 -420 1006 -416
rect 1139 -424 1143 -420
rect 1147 -423 1151 -419
rect 1428 -422 1432 -416
rect 1436 -422 1440 -416
rect 1893 -426 1897 -422
rect 1901 -425 1905 -421
rect 1992 -423 1996 -419
rect 2000 -422 2004 -418
rect 2098 -420 2102 -416
rect 2106 -419 2110 -415
rect 611 -449 615 -443
rect 619 -449 623 -443
rect 1602 -447 1606 -438
rect 1610 -447 1614 -438
rect 1843 -439 1847 -430
rect 1851 -439 1855 -430
rect 1957 -440 1961 -434
rect 1965 -440 1969 -434
rect 1939 -447 1943 -441
rect 1947 -447 1951 -441
rect 2069 -440 2073 -434
rect 2077 -440 2081 -434
rect 2051 -447 2055 -441
rect 2059 -447 2063 -441
rect 1722 -454 1726 -448
rect 1730 -454 1734 -448
rect 1759 -452 1763 -448
rect 1767 -451 1771 -447
rect 1602 -467 1606 -458
rect 1610 -467 1614 -458
rect 1843 -459 1847 -450
rect 1851 -459 1855 -450
rect 1699 -467 1703 -461
rect 1707 -467 1711 -461
rect 689 -480 693 -474
rect 697 -480 701 -474
rect 1722 -480 1726 -474
rect 1730 -480 1734 -474
rect 1602 -495 1606 -486
rect 1610 -495 1614 -486
rect 1843 -487 1847 -478
rect 1851 -487 1855 -478
rect 689 -506 693 -500
rect 697 -506 701 -500
rect 1007 -506 1011 -500
rect 1015 -506 1019 -500
rect 1044 -523 1048 -519
rect 1052 -522 1056 -518
rect 1602 -515 1606 -506
rect 1610 -515 1614 -506
rect 1139 -526 1143 -520
rect 1147 -526 1151 -520
rect 1176 -524 1180 -520
rect 1184 -523 1188 -519
rect 1007 -532 1011 -526
rect 1015 -532 1019 -526
rect 1116 -539 1120 -533
rect 1124 -539 1128 -533
rect 1653 -538 1657 -534
rect 1661 -537 1665 -533
rect 1139 -552 1143 -546
rect 1147 -552 1151 -546
rect 612 -559 616 -553
rect 620 -559 624 -553
rect 612 -585 616 -579
rect 620 -585 624 -579
rect 1101 -706 1105 -700
rect 1118 -706 1122 -700
rect 1046 -718 1050 -714
rect 1054 -717 1058 -713
rect 1361 -709 1365 -703
rect 1378 -709 1382 -703
rect 1306 -721 1310 -717
rect 1314 -720 1318 -716
rect 1135 -735 1139 -731
rect 1143 -734 1147 -730
rect 1395 -738 1399 -734
rect 1403 -737 1407 -733
rect 1101 -747 1106 -741
rect 1118 -747 1122 -741
rect 1361 -750 1366 -744
rect 1378 -750 1382 -744
rect 1046 -770 1050 -766
rect 1054 -769 1058 -765
rect 1306 -773 1310 -769
rect 1314 -772 1318 -768
rect 1059 -849 1063 -843
rect 1067 -849 1071 -843
rect 1096 -866 1100 -862
rect 1104 -865 1108 -861
rect 1059 -875 1063 -869
rect 1067 -875 1071 -869
rect 1370 -873 1374 -864
rect 1378 -873 1382 -864
rect 1462 -874 1466 -868
rect 1470 -874 1474 -868
rect 1444 -881 1448 -875
rect 1452 -881 1456 -875
rect 1215 -888 1219 -882
rect 1223 -888 1227 -882
rect 1252 -886 1256 -882
rect 1260 -885 1264 -881
rect 1370 -893 1374 -884
rect 1378 -893 1382 -884
rect 1192 -901 1196 -895
rect 1200 -901 1204 -895
rect 1215 -914 1219 -908
rect 1223 -914 1227 -908
rect 1370 -921 1374 -912
rect 1378 -921 1382 -912
<< pdcontact >>
rect 1415 -241 1419 -235
rect 1423 -241 1427 -235
rect 1675 -244 1679 -238
rect 1683 -244 1687 -238
rect 1504 -258 1508 -252
rect 1512 -258 1516 -252
rect 1764 -261 1768 -255
rect 1772 -261 1776 -255
rect 488 -287 492 -281
rect 496 -287 500 -281
rect 657 -290 661 -284
rect 665 -290 669 -284
rect 577 -304 581 -298
rect 585 -304 589 -298
rect 1415 -293 1419 -287
rect 1423 -293 1427 -287
rect 1675 -296 1679 -290
rect 1683 -296 1687 -290
rect 722 -307 726 -301
rect 730 -307 734 -301
rect 488 -339 492 -333
rect 496 -339 500 -333
rect 657 -342 661 -336
rect 665 -342 669 -336
rect 994 -351 998 -345
rect 1002 -351 1006 -345
rect 1420 -347 1424 -341
rect 1428 -347 1432 -341
rect 1139 -354 1143 -348
rect 1147 -354 1151 -348
rect 603 -374 607 -368
rect 611 -374 615 -368
rect 1069 -368 1073 -362
rect 1077 -368 1081 -362
rect 1446 -363 1450 -357
rect 1454 -363 1458 -357
rect 1635 -361 1639 -349
rect 1643 -361 1647 -349
rect 1228 -371 1232 -365
rect 1236 -371 1240 -365
rect 629 -390 633 -384
rect 637 -390 641 -384
rect 1618 -381 1622 -369
rect 1626 -381 1630 -369
rect 994 -403 998 -397
rect 1002 -403 1006 -397
rect 1139 -406 1143 -400
rect 1147 -406 1151 -400
rect 1465 -395 1469 -389
rect 1473 -395 1477 -389
rect 1598 -395 1602 -383
rect 1606 -395 1610 -383
rect 1706 -385 1710 -373
rect 1714 -385 1718 -373
rect 1859 -373 1863 -361
rect 1867 -373 1871 -361
rect 1839 -387 1843 -375
rect 1847 -387 1851 -375
rect 1947 -384 1951 -372
rect 1955 -384 1959 -372
rect 2059 -384 2063 -372
rect 2067 -384 2071 -372
rect 1579 -413 1583 -401
rect 1587 -413 1591 -401
rect 1820 -405 1824 -393
rect 1828 -405 1832 -393
rect 1698 -419 1702 -407
rect 1706 -419 1710 -407
rect 1729 -419 1733 -407
rect 1737 -419 1741 -407
rect 1893 -408 1897 -402
rect 1901 -408 1905 -402
rect 681 -431 685 -425
rect 689 -431 693 -425
rect 1947 -416 1951 -404
rect 1955 -416 1959 -404
rect 1992 -405 1996 -399
rect 2000 -405 2004 -399
rect 2098 -402 2102 -396
rect 2106 -402 2110 -396
rect 2059 -416 2063 -404
rect 2067 -416 2071 -404
rect 1759 -434 1763 -428
rect 1767 -434 1771 -428
rect 707 -447 711 -441
rect 715 -447 719 -441
rect 999 -457 1003 -451
rect 1007 -457 1011 -451
rect 1123 -457 1127 -445
rect 1131 -457 1135 -445
rect 1025 -473 1029 -467
rect 1033 -473 1037 -467
rect 1115 -491 1119 -479
rect 1123 -491 1127 -479
rect 1146 -491 1150 -479
rect 1154 -491 1158 -479
rect 604 -510 608 -504
rect 612 -510 616 -504
rect 1044 -505 1048 -499
rect 1052 -505 1056 -499
rect 1176 -506 1180 -500
rect 1184 -506 1188 -500
rect 630 -526 634 -520
rect 638 -526 642 -520
rect 1653 -520 1657 -514
rect 1661 -520 1665 -514
rect 1046 -700 1050 -694
rect 1054 -700 1058 -694
rect 1306 -703 1310 -697
rect 1314 -703 1318 -697
rect 1135 -717 1139 -711
rect 1143 -717 1147 -711
rect 1395 -720 1399 -714
rect 1403 -720 1407 -714
rect 1046 -752 1050 -746
rect 1054 -752 1058 -746
rect 1306 -755 1310 -749
rect 1314 -755 1318 -749
rect 1051 -800 1055 -794
rect 1059 -800 1063 -794
rect 1077 -816 1081 -810
rect 1085 -816 1089 -810
rect 1199 -819 1203 -807
rect 1207 -819 1211 -807
rect 1386 -807 1390 -795
rect 1394 -807 1398 -795
rect 1366 -821 1370 -809
rect 1374 -821 1378 -809
rect 1452 -818 1456 -806
rect 1460 -818 1464 -806
rect 1347 -839 1351 -827
rect 1355 -839 1359 -827
rect 1096 -848 1100 -842
rect 1104 -848 1108 -842
rect 1191 -853 1195 -841
rect 1199 -853 1203 -841
rect 1222 -853 1226 -841
rect 1230 -853 1234 -841
rect 1452 -850 1456 -838
rect 1460 -850 1464 -838
rect 1252 -868 1256 -862
rect 1260 -868 1264 -862
<< polysilicon >>
rect 1420 -235 1422 -232
rect 1680 -238 1682 -235
rect 1479 -241 1481 -238
rect 1420 -255 1422 -241
rect 1739 -244 1741 -241
rect 1479 -256 1481 -247
rect 1509 -252 1511 -249
rect 1680 -258 1682 -244
rect 1420 -261 1422 -258
rect 1509 -272 1511 -258
rect 1739 -259 1741 -250
rect 1769 -255 1771 -252
rect 1680 -264 1682 -261
rect 1769 -275 1771 -261
rect 1509 -278 1511 -275
rect 493 -281 495 -278
rect 662 -284 664 -281
rect 1479 -282 1481 -279
rect 1769 -281 1771 -278
rect 552 -287 554 -284
rect 493 -301 495 -287
rect 1420 -287 1422 -284
rect 697 -290 699 -287
rect 552 -302 554 -293
rect 582 -298 584 -295
rect 662 -304 664 -290
rect 1739 -285 1741 -282
rect 493 -307 495 -304
rect 582 -318 584 -304
rect 697 -305 699 -296
rect 727 -301 729 -298
rect 1420 -300 1422 -293
rect 1479 -297 1481 -288
rect 1680 -290 1682 -287
rect 1419 -304 1422 -300
rect 1680 -303 1682 -296
rect 1739 -300 1741 -291
rect 1420 -307 1422 -304
rect 662 -310 664 -307
rect 727 -321 729 -307
rect 1679 -307 1682 -303
rect 1680 -310 1682 -307
rect 1420 -313 1422 -310
rect 1680 -316 1682 -313
rect 582 -324 584 -321
rect 552 -328 554 -325
rect 727 -327 729 -324
rect 493 -333 495 -330
rect 697 -331 699 -328
rect 493 -346 495 -339
rect 552 -343 554 -334
rect 662 -336 664 -333
rect 492 -350 495 -346
rect 662 -349 664 -342
rect 697 -346 699 -337
rect 1425 -341 1427 -338
rect 999 -345 1001 -342
rect 493 -353 495 -350
rect 661 -353 664 -349
rect 1144 -348 1146 -345
rect 1044 -351 1046 -348
rect 662 -356 664 -353
rect 493 -359 495 -356
rect 662 -362 664 -359
rect 999 -365 1001 -351
rect 1203 -354 1205 -351
rect 1425 -354 1427 -347
rect 1640 -349 1642 -342
rect 608 -368 610 -365
rect 1044 -366 1046 -357
rect 1074 -362 1076 -359
rect 1144 -368 1146 -354
rect 1451 -357 1453 -350
rect 999 -371 1001 -368
rect 608 -381 610 -374
rect 634 -384 636 -377
rect 1074 -382 1076 -368
rect 1203 -369 1205 -360
rect 1233 -365 1235 -362
rect 1864 -361 1866 -354
rect 1451 -366 1453 -363
rect 1623 -369 1625 -362
rect 1640 -364 1642 -361
rect 1144 -374 1146 -371
rect 1233 -385 1235 -371
rect 1603 -383 1605 -376
rect 1711 -373 1713 -366
rect 1074 -388 1076 -385
rect 634 -393 636 -390
rect 1044 -392 1046 -389
rect 1233 -391 1235 -388
rect 1433 -390 1435 -383
rect 1470 -389 1472 -386
rect 999 -397 1001 -394
rect 1203 -395 1205 -392
rect 999 -410 1001 -403
rect 1044 -407 1046 -398
rect 1144 -400 1146 -397
rect 1433 -399 1435 -396
rect 616 -417 618 -410
rect 998 -414 1001 -410
rect 1144 -413 1146 -406
rect 1203 -410 1205 -401
rect 1470 -409 1472 -395
rect 1584 -401 1586 -394
rect 1623 -384 1625 -381
rect 1844 -375 1846 -368
rect 1952 -372 1954 -365
rect 2064 -372 2066 -365
rect 1711 -388 1713 -385
rect 1825 -393 1827 -386
rect 1864 -376 1866 -373
rect 1952 -387 1954 -384
rect 2064 -387 2066 -384
rect 1844 -390 1846 -387
rect 1603 -398 1605 -395
rect 999 -417 1001 -414
rect 1143 -417 1146 -413
rect 1433 -416 1435 -413
rect 1470 -415 1472 -412
rect 1703 -407 1705 -400
rect 1734 -407 1736 -404
rect 2103 -396 2105 -393
rect 1898 -402 1900 -399
rect 1584 -416 1586 -413
rect 1144 -420 1146 -417
rect 616 -426 618 -423
rect 686 -425 688 -422
rect 999 -423 1001 -420
rect 1825 -408 1827 -405
rect 1952 -404 1954 -397
rect 1997 -399 1999 -396
rect 1703 -422 1705 -419
rect 1144 -426 1146 -423
rect 1433 -429 1435 -422
rect 1734 -426 1736 -419
rect 1898 -422 1900 -408
rect 2064 -404 2066 -397
rect 1952 -419 1954 -416
rect 1997 -419 1999 -405
rect 2103 -416 2105 -402
rect 1764 -428 1766 -425
rect 686 -438 688 -431
rect 616 -443 618 -440
rect 712 -441 714 -434
rect 1607 -438 1609 -431
rect 1848 -430 1850 -423
rect 2064 -419 2066 -416
rect 2103 -422 2105 -419
rect 1997 -425 1999 -422
rect 1898 -428 1900 -425
rect 1128 -445 1130 -438
rect 616 -456 618 -449
rect 712 -450 714 -447
rect 1004 -451 1006 -448
rect 1607 -450 1609 -447
rect 1727 -448 1729 -441
rect 1764 -448 1766 -434
rect 1962 -434 1964 -431
rect 2074 -434 2076 -431
rect 1848 -442 1850 -439
rect 1944 -441 1946 -434
rect 1962 -447 1964 -440
rect 2056 -441 2058 -434
rect 2074 -447 2076 -440
rect 1848 -450 1850 -447
rect 1944 -450 1946 -447
rect 2056 -450 2058 -447
rect 1764 -454 1766 -451
rect 1004 -464 1006 -457
rect 1128 -460 1130 -457
rect 1607 -458 1609 -455
rect 1727 -457 1729 -454
rect 1030 -467 1032 -460
rect 1704 -461 1706 -458
rect 1848 -466 1850 -459
rect 694 -474 696 -467
rect 1030 -476 1032 -473
rect 1120 -479 1122 -472
rect 1607 -474 1609 -467
rect 1704 -474 1706 -467
rect 1727 -474 1729 -471
rect 1151 -479 1153 -476
rect 694 -483 696 -480
rect 1607 -486 1609 -479
rect 1848 -478 1850 -471
rect 694 -500 696 -497
rect 1012 -500 1014 -493
rect 1120 -494 1122 -491
rect 1049 -499 1051 -496
rect 1151 -498 1153 -491
rect 1727 -487 1729 -480
rect 1848 -490 1850 -487
rect 609 -504 611 -501
rect 1181 -500 1183 -497
rect 1607 -498 1609 -495
rect 609 -517 611 -510
rect 694 -513 696 -506
rect 1012 -509 1014 -506
rect 635 -520 637 -513
rect 1049 -519 1051 -505
rect 1607 -506 1609 -503
rect 1144 -520 1146 -513
rect 1181 -520 1183 -506
rect 1658 -514 1660 -511
rect 1012 -526 1014 -523
rect 1049 -525 1051 -522
rect 1607 -522 1609 -515
rect 1181 -526 1183 -523
rect 635 -529 637 -526
rect 1144 -529 1146 -526
rect 1012 -539 1014 -532
rect 1121 -533 1123 -530
rect 1658 -534 1660 -520
rect 1121 -546 1123 -539
rect 1658 -540 1660 -537
rect 1144 -546 1146 -543
rect 617 -553 619 -546
rect 1144 -559 1146 -552
rect 617 -562 619 -559
rect 617 -579 619 -576
rect 617 -592 619 -585
rect 1051 -694 1053 -691
rect 1311 -697 1313 -694
rect 1110 -700 1112 -697
rect 1051 -714 1053 -700
rect 1370 -703 1372 -700
rect 1110 -715 1112 -706
rect 1140 -711 1142 -708
rect 1311 -717 1313 -703
rect 1051 -720 1053 -717
rect 1140 -731 1142 -717
rect 1370 -718 1372 -709
rect 1400 -714 1402 -711
rect 1311 -723 1313 -720
rect 1400 -734 1402 -720
rect 1140 -737 1142 -734
rect 1110 -741 1112 -738
rect 1400 -740 1402 -737
rect 1051 -746 1053 -743
rect 1370 -744 1372 -741
rect 1051 -759 1053 -752
rect 1110 -756 1112 -747
rect 1311 -749 1313 -746
rect 1050 -763 1053 -759
rect 1311 -762 1313 -755
rect 1370 -759 1372 -750
rect 1051 -766 1053 -763
rect 1310 -766 1313 -762
rect 1311 -769 1313 -766
rect 1051 -772 1053 -769
rect 1311 -775 1313 -772
rect 1056 -794 1058 -791
rect 1391 -795 1393 -788
rect 1056 -807 1058 -800
rect 1082 -810 1084 -803
rect 1204 -807 1206 -800
rect 1082 -819 1084 -816
rect 1371 -809 1373 -802
rect 1457 -806 1459 -799
rect 1204 -822 1206 -819
rect 1352 -827 1354 -820
rect 1391 -810 1393 -807
rect 1457 -821 1459 -818
rect 1371 -824 1373 -821
rect 1064 -843 1066 -836
rect 1101 -842 1103 -839
rect 1196 -841 1198 -834
rect 1227 -841 1229 -838
rect 1457 -838 1459 -831
rect 1064 -852 1066 -849
rect 1101 -862 1103 -848
rect 1352 -842 1354 -839
rect 1457 -853 1459 -850
rect 1196 -856 1198 -853
rect 1227 -860 1229 -853
rect 1257 -862 1259 -859
rect 1064 -869 1066 -866
rect 1101 -868 1103 -865
rect 1375 -864 1377 -857
rect 1064 -882 1066 -875
rect 1220 -882 1222 -875
rect 1257 -882 1259 -868
rect 1467 -868 1469 -865
rect 1375 -876 1377 -873
rect 1449 -875 1451 -868
rect 1467 -881 1469 -874
rect 1375 -884 1377 -881
rect 1449 -884 1451 -881
rect 1257 -888 1259 -885
rect 1220 -891 1222 -888
rect 1197 -895 1199 -892
rect 1375 -900 1377 -893
rect 1197 -908 1199 -901
rect 1220 -908 1222 -905
rect 1375 -912 1377 -905
rect 1220 -921 1222 -914
rect 1375 -924 1377 -921
<< polycontact >>
rect 1416 -252 1420 -248
rect 1475 -256 1479 -251
rect 1676 -255 1680 -251
rect 1505 -269 1509 -265
rect 1735 -259 1739 -254
rect 1765 -272 1769 -268
rect 489 -298 493 -294
rect 548 -302 552 -297
rect 658 -301 662 -297
rect 578 -315 582 -311
rect 693 -305 697 -300
rect 1475 -297 1479 -293
rect 1415 -304 1419 -300
rect 1735 -300 1739 -296
rect 723 -318 727 -314
rect 1675 -307 1679 -303
rect 548 -343 552 -339
rect 488 -350 492 -346
rect 693 -346 697 -342
rect 657 -353 661 -349
rect 1636 -346 1640 -342
rect 995 -362 999 -358
rect 1421 -354 1425 -350
rect 1447 -354 1451 -350
rect 1040 -366 1044 -361
rect 1140 -365 1144 -361
rect 604 -381 608 -377
rect 630 -381 634 -377
rect 1070 -379 1074 -375
rect 1199 -369 1203 -364
rect 1860 -358 1864 -354
rect 1619 -366 1623 -362
rect 1229 -382 1233 -378
rect 1599 -380 1603 -376
rect 1707 -370 1711 -366
rect 1840 -372 1844 -368
rect 1429 -387 1433 -383
rect 1040 -407 1044 -403
rect 612 -414 616 -410
rect 994 -414 998 -410
rect 1199 -410 1203 -406
rect 1466 -406 1470 -402
rect 1580 -398 1584 -394
rect 1948 -369 1952 -365
rect 2060 -369 2064 -365
rect 1821 -390 1825 -386
rect 1139 -417 1143 -413
rect 1699 -404 1703 -400
rect 1948 -401 1952 -397
rect 1894 -419 1898 -415
rect 1429 -429 1433 -425
rect 1730 -426 1734 -422
rect 2060 -401 2064 -397
rect 1993 -416 1997 -412
rect 2099 -413 2103 -409
rect 1844 -427 1848 -423
rect 682 -438 686 -434
rect 708 -438 712 -434
rect 1603 -435 1607 -431
rect 1124 -442 1128 -438
rect 612 -456 616 -452
rect 1723 -445 1727 -441
rect 1760 -445 1764 -441
rect 1940 -438 1944 -434
rect 2052 -438 2056 -434
rect 1958 -447 1962 -443
rect 2070 -447 2074 -443
rect 1000 -464 1004 -460
rect 1026 -464 1030 -460
rect 1844 -466 1848 -462
rect 690 -471 694 -467
rect 1116 -476 1120 -472
rect 1603 -474 1607 -470
rect 1700 -474 1704 -470
rect 1603 -483 1607 -479
rect 1844 -475 1848 -471
rect 1008 -497 1012 -493
rect 1147 -498 1151 -494
rect 1723 -487 1727 -483
rect 605 -517 609 -513
rect 690 -513 694 -509
rect 631 -517 635 -513
rect 1045 -516 1049 -512
rect 1140 -517 1144 -513
rect 1177 -517 1181 -513
rect 1603 -522 1607 -518
rect 1008 -539 1012 -535
rect 1654 -531 1658 -527
rect 1117 -546 1121 -542
rect 613 -550 617 -546
rect 1140 -559 1144 -555
rect 613 -592 617 -588
rect 1047 -711 1051 -707
rect 1106 -715 1110 -710
rect 1307 -714 1311 -710
rect 1136 -728 1140 -724
rect 1366 -718 1370 -713
rect 1396 -731 1400 -727
rect 1106 -756 1110 -752
rect 1046 -763 1050 -759
rect 1366 -759 1370 -755
rect 1306 -766 1310 -762
rect 1387 -792 1391 -788
rect 1052 -807 1056 -803
rect 1078 -807 1082 -803
rect 1200 -804 1204 -800
rect 1367 -806 1371 -802
rect 1453 -803 1457 -799
rect 1348 -824 1352 -820
rect 1060 -840 1064 -836
rect 1192 -838 1196 -834
rect 1453 -835 1457 -831
rect 1097 -859 1101 -855
rect 1223 -860 1227 -856
rect 1371 -861 1375 -857
rect 1060 -882 1064 -878
rect 1216 -879 1220 -875
rect 1253 -879 1257 -875
rect 1445 -872 1449 -868
rect 1463 -881 1467 -877
rect 1371 -900 1375 -896
rect 1193 -908 1197 -904
rect 1371 -909 1375 -905
rect 1216 -921 1220 -917
<< metal1 >>
rect 1400 -221 1474 -216
rect 1400 -248 1404 -221
rect 1409 -230 1433 -226
rect 1415 -235 1419 -230
rect 1470 -241 1474 -221
rect 1660 -224 1734 -219
rect 1498 -247 1522 -243
rect 1380 -252 1416 -248
rect 473 -267 547 -262
rect 473 -294 477 -267
rect 482 -276 506 -272
rect 488 -281 492 -276
rect 543 -287 547 -267
rect 642 -270 692 -265
rect 571 -293 595 -289
rect 453 -298 489 -294
rect 488 -308 492 -305
rect 482 -312 506 -308
rect 560 -311 564 -293
rect 577 -298 581 -293
rect 642 -297 646 -270
rect 651 -279 675 -275
rect 657 -284 661 -279
rect 688 -290 692 -270
rect 716 -296 740 -292
rect 585 -310 589 -304
rect 642 -301 658 -297
rect 642 -310 646 -301
rect 560 -315 578 -311
rect 585 -314 646 -310
rect 657 -311 661 -308
rect 482 -328 506 -324
rect 560 -328 564 -315
rect 585 -317 589 -314
rect 577 -325 581 -322
rect 488 -333 492 -328
rect 571 -329 595 -325
rect 488 -360 492 -357
rect 619 -358 623 -314
rect 651 -315 675 -311
rect 705 -314 709 -296
rect 722 -301 726 -296
rect 705 -318 723 -314
rect 651 -331 675 -327
rect 705 -331 709 -318
rect 722 -328 726 -325
rect 657 -336 661 -331
rect 716 -332 740 -328
rect 979 -331 1039 -326
rect 482 -364 506 -360
rect 576 -362 623 -358
rect 576 -452 580 -362
rect 587 -381 604 -377
rect 587 -409 591 -381
rect 611 -398 615 -374
rect 619 -377 623 -362
rect 979 -358 983 -331
rect 988 -340 1012 -336
rect 994 -345 998 -340
rect 1035 -351 1039 -331
rect 1124 -334 1198 -329
rect 1063 -357 1087 -353
rect 657 -363 661 -360
rect 959 -362 995 -358
rect 651 -367 675 -363
rect 619 -381 630 -377
rect 637 -398 641 -390
rect 611 -402 641 -398
rect 592 -414 612 -410
rect 619 -417 623 -402
rect 654 -419 701 -415
rect 611 -443 615 -423
rect 562 -456 612 -452
rect 577 -498 624 -494
rect 577 -588 581 -498
rect 588 -517 605 -513
rect 588 -545 592 -517
rect 612 -534 616 -510
rect 620 -513 624 -498
rect 654 -509 658 -419
rect 665 -438 682 -434
rect 665 -466 669 -438
rect 689 -455 693 -431
rect 697 -434 701 -419
rect 697 -438 708 -434
rect 972 -441 976 -362
rect 994 -372 998 -369
rect 988 -376 1012 -372
rect 1052 -375 1056 -357
rect 1069 -362 1073 -357
rect 1124 -361 1128 -334
rect 1133 -343 1157 -339
rect 1139 -348 1143 -343
rect 1194 -354 1198 -334
rect 1393 -331 1397 -252
rect 1415 -262 1419 -259
rect 1409 -266 1433 -262
rect 1487 -265 1491 -247
rect 1504 -252 1508 -247
rect 1660 -251 1664 -224
rect 1669 -233 1693 -229
rect 1675 -238 1679 -233
rect 1730 -244 1734 -224
rect 1758 -250 1782 -246
rect 1512 -264 1516 -258
rect 1639 -255 1676 -251
rect 1639 -264 1643 -255
rect 1487 -269 1505 -265
rect 1512 -268 1643 -264
rect 1675 -265 1679 -262
rect 1409 -282 1433 -278
rect 1487 -282 1491 -269
rect 1512 -271 1516 -268
rect 1504 -279 1508 -276
rect 1415 -287 1419 -282
rect 1498 -283 1522 -279
rect 1415 -314 1419 -311
rect 1409 -318 1433 -314
rect 1393 -335 1440 -331
rect 1222 -360 1246 -356
rect 1077 -374 1081 -368
rect 1103 -365 1140 -361
rect 1103 -374 1107 -365
rect 1052 -379 1070 -375
rect 1077 -378 1096 -374
rect 988 -392 1012 -388
rect 1052 -392 1056 -379
rect 1077 -381 1081 -378
rect 1101 -378 1107 -374
rect 1139 -375 1143 -372
rect 1133 -379 1157 -375
rect 1211 -378 1215 -360
rect 1228 -365 1232 -360
rect 1211 -382 1229 -378
rect 1069 -389 1073 -386
rect 994 -397 998 -392
rect 1063 -393 1087 -389
rect 1133 -395 1157 -391
rect 1211 -395 1215 -382
rect 1228 -392 1232 -389
rect 1139 -400 1143 -395
rect 1222 -396 1246 -392
rect 994 -424 998 -421
rect 988 -428 1012 -424
rect 1139 -427 1143 -424
rect 1393 -425 1397 -335
rect 1404 -354 1421 -350
rect 1404 -382 1408 -354
rect 1428 -371 1432 -347
rect 1436 -350 1440 -335
rect 1557 -342 1561 -268
rect 1669 -269 1693 -265
rect 1747 -268 1751 -250
rect 1764 -255 1768 -250
rect 1747 -272 1765 -268
rect 1669 -285 1693 -281
rect 1747 -285 1751 -272
rect 1764 -282 1768 -279
rect 1675 -290 1679 -285
rect 1758 -286 1782 -282
rect 1675 -317 1679 -314
rect 1669 -321 1693 -317
rect 1538 -346 1636 -342
rect 1436 -354 1447 -350
rect 1454 -371 1458 -363
rect 1428 -375 1458 -371
rect 1409 -387 1429 -383
rect 1436 -390 1440 -375
rect 1428 -416 1432 -396
rect 1449 -402 1453 -375
rect 1459 -384 1483 -380
rect 1465 -389 1469 -384
rect 1473 -402 1477 -395
rect 1449 -406 1466 -402
rect 1473 -406 1485 -402
rect 1473 -408 1477 -406
rect 1465 -416 1469 -413
rect 1459 -420 1483 -416
rect 1133 -431 1157 -427
rect 1393 -429 1429 -425
rect 715 -455 719 -447
rect 689 -459 719 -455
rect 972 -445 1019 -441
rect 670 -471 690 -467
rect 697 -474 701 -459
rect 689 -500 693 -480
rect 654 -513 690 -509
rect 620 -517 631 -513
rect 638 -534 642 -526
rect 654 -534 657 -513
rect 612 -538 657 -534
rect 972 -535 976 -445
rect 983 -464 1000 -460
rect 983 -492 987 -464
rect 1007 -481 1011 -457
rect 1015 -460 1019 -445
rect 1084 -442 1124 -438
rect 1015 -464 1026 -460
rect 1033 -481 1037 -473
rect 1007 -485 1037 -481
rect 988 -497 1008 -493
rect 1015 -500 1019 -485
rect 1007 -526 1011 -506
rect 1028 -512 1032 -485
rect 1038 -494 1062 -490
rect 1044 -499 1048 -494
rect 1052 -512 1056 -505
rect 1084 -512 1088 -442
rect 1123 -469 1127 -457
rect 1123 -473 1150 -469
rect 1123 -479 1127 -473
rect 1146 -479 1150 -473
rect 1115 -504 1119 -491
rect 1154 -504 1158 -491
rect 1170 -495 1194 -491
rect 1115 -508 1158 -504
rect 1176 -500 1180 -495
rect 1028 -516 1045 -512
rect 1052 -516 1088 -512
rect 1052 -518 1056 -516
rect 1044 -526 1048 -523
rect 1038 -530 1062 -526
rect 593 -550 613 -546
rect 620 -553 624 -538
rect 972 -539 1008 -535
rect 1084 -542 1088 -516
rect 1116 -533 1120 -508
rect 1147 -520 1151 -508
rect 1154 -513 1158 -508
rect 1154 -517 1177 -513
rect 1538 -518 1542 -346
rect 1550 -366 1619 -362
rect 1550 -479 1554 -366
rect 1561 -380 1599 -376
rect 1561 -470 1565 -380
rect 1571 -398 1580 -394
rect 1571 -431 1575 -398
rect 1587 -423 1591 -413
rect 1606 -423 1610 -395
rect 1626 -423 1630 -381
rect 1643 -423 1647 -361
rect 1791 -358 1860 -354
rect 1587 -427 1647 -423
rect 1667 -370 1707 -366
rect 1571 -435 1603 -431
rect 1610 -438 1614 -427
rect 1602 -458 1606 -447
rect 1561 -474 1603 -470
rect 1550 -483 1603 -479
rect 1610 -486 1614 -467
rect 1602 -506 1606 -495
rect 1538 -522 1603 -518
rect 1084 -546 1117 -542
rect 1139 -546 1143 -526
rect 1176 -527 1180 -524
rect 1639 -527 1643 -427
rect 1667 -470 1671 -370
rect 1706 -397 1710 -385
rect 1706 -401 1733 -397
rect 1706 -407 1710 -401
rect 1729 -407 1733 -401
rect 1698 -432 1702 -419
rect 1737 -432 1741 -419
rect 1753 -423 1777 -419
rect 1698 -436 1741 -432
rect 1759 -428 1763 -423
rect 1699 -461 1703 -436
rect 1730 -448 1734 -436
rect 1737 -441 1741 -436
rect 1737 -445 1760 -441
rect 1667 -474 1700 -470
rect 1722 -474 1726 -454
rect 1759 -455 1763 -452
rect 1753 -459 1777 -455
rect 1791 -471 1795 -358
rect 1802 -372 1840 -368
rect 1802 -462 1806 -372
rect 1812 -390 1821 -386
rect 1812 -423 1816 -390
rect 1828 -415 1832 -405
rect 1847 -415 1851 -387
rect 1867 -415 1871 -373
rect 1915 -369 1948 -365
rect 2023 -369 2060 -365
rect 1887 -397 1911 -393
rect 1893 -402 1897 -397
rect 1901 -415 1905 -408
rect 1915 -415 1919 -369
rect 1927 -401 1948 -397
rect 1955 -404 1959 -384
rect 1986 -394 2010 -390
rect 1828 -419 1894 -415
rect 1901 -419 1919 -415
rect 1812 -427 1844 -423
rect 1851 -430 1855 -419
rect 1901 -421 1905 -419
rect 1893 -429 1897 -426
rect 1887 -433 1911 -429
rect 1843 -450 1847 -439
rect 1915 -450 1919 -419
rect 1992 -399 1996 -394
rect 2000 -412 2004 -405
rect 2023 -412 2027 -369
rect 1973 -416 1993 -412
rect 2000 -416 2027 -412
rect 1947 -424 1951 -416
rect 1973 -424 1976 -416
rect 2000 -418 2004 -416
rect 1947 -428 1976 -424
rect 1992 -426 1996 -423
rect 2023 -424 2027 -416
rect 2035 -401 2060 -397
rect 1927 -438 1940 -434
rect 1947 -441 1951 -428
rect 1957 -434 1961 -428
rect 1986 -430 2010 -426
rect 2023 -428 2030 -424
rect 2026 -433 2030 -428
rect 1958 -450 1962 -447
rect 1915 -454 1962 -450
rect 2035 -450 2040 -401
rect 2067 -404 2071 -384
rect 2092 -391 2116 -387
rect 2098 -396 2102 -391
rect 2080 -413 2099 -409
rect 2059 -424 2063 -416
rect 2080 -424 2084 -413
rect 2098 -423 2102 -420
rect 2059 -428 2084 -424
rect 2092 -427 2116 -423
rect 2059 -441 2063 -428
rect 2069 -434 2073 -428
rect 2070 -450 2074 -447
rect 2035 -454 2074 -450
rect 1802 -466 1844 -462
rect 1791 -475 1844 -471
rect 1851 -478 1855 -459
rect 1647 -509 1671 -505
rect 1653 -514 1657 -509
rect 1661 -527 1665 -520
rect 2035 -527 2040 -454
rect 1170 -531 1194 -527
rect 1639 -531 1654 -527
rect 1661 -531 2040 -527
rect 1661 -533 1665 -531
rect 1653 -540 1657 -538
rect 612 -579 616 -559
rect 563 -592 613 -588
rect 1031 -680 1105 -675
rect 1031 -707 1035 -680
rect 1040 -689 1064 -685
rect 1046 -694 1050 -689
rect 1101 -700 1105 -680
rect 1291 -683 1365 -678
rect 1129 -706 1153 -702
rect 1011 -711 1047 -707
rect 1024 -784 1028 -711
rect 1046 -721 1050 -718
rect 1040 -725 1064 -721
rect 1118 -724 1122 -706
rect 1135 -711 1139 -706
rect 1291 -710 1295 -683
rect 1300 -692 1324 -688
rect 1306 -697 1310 -692
rect 1361 -703 1365 -683
rect 1389 -709 1413 -705
rect 1143 -723 1147 -717
rect 1270 -714 1307 -710
rect 1270 -723 1274 -714
rect 1118 -728 1136 -724
rect 1143 -727 1171 -723
rect 1040 -741 1064 -737
rect 1118 -741 1122 -728
rect 1143 -730 1147 -727
rect 1176 -727 1274 -723
rect 1306 -724 1310 -721
rect 1135 -738 1139 -735
rect 1046 -746 1050 -741
rect 1129 -742 1153 -738
rect 1046 -773 1050 -770
rect 1040 -777 1064 -773
rect 1024 -788 1071 -784
rect 1024 -878 1028 -788
rect 1035 -807 1052 -803
rect 1035 -835 1039 -807
rect 1059 -824 1063 -800
rect 1067 -803 1071 -788
rect 1261 -788 1265 -727
rect 1300 -728 1324 -724
rect 1378 -727 1382 -709
rect 1395 -714 1399 -709
rect 1378 -731 1396 -727
rect 1300 -744 1324 -740
rect 1378 -744 1382 -731
rect 1395 -741 1399 -738
rect 1306 -749 1310 -744
rect 1389 -745 1413 -741
rect 1306 -776 1310 -773
rect 1300 -780 1324 -776
rect 1261 -792 1387 -788
rect 1067 -807 1078 -803
rect 1160 -804 1200 -800
rect 1160 -808 1164 -804
rect 1085 -824 1089 -816
rect 1059 -828 1089 -824
rect 1128 -812 1164 -808
rect 1040 -840 1060 -836
rect 1067 -843 1071 -828
rect 1059 -869 1063 -849
rect 1080 -855 1084 -828
rect 1090 -837 1114 -833
rect 1096 -842 1100 -837
rect 1104 -855 1108 -848
rect 1128 -855 1132 -812
rect 1080 -859 1097 -855
rect 1104 -859 1132 -855
rect 1104 -861 1108 -859
rect 1096 -869 1100 -866
rect 1090 -873 1114 -869
rect 1024 -882 1060 -878
rect 1160 -904 1164 -812
rect 1199 -831 1203 -819
rect 1199 -835 1226 -831
rect 1199 -841 1203 -835
rect 1222 -841 1226 -835
rect 1191 -866 1195 -853
rect 1230 -866 1234 -853
rect 1246 -857 1270 -853
rect 1191 -870 1234 -866
rect 1252 -862 1256 -857
rect 1192 -895 1196 -870
rect 1223 -882 1227 -870
rect 1230 -875 1234 -870
rect 1230 -879 1253 -875
rect 1160 -908 1193 -904
rect 1215 -908 1219 -888
rect 1252 -889 1256 -886
rect 1246 -893 1270 -889
rect 1318 -905 1322 -792
rect 1329 -806 1367 -802
rect 1329 -896 1333 -806
rect 1339 -824 1348 -820
rect 1339 -857 1343 -824
rect 1355 -849 1359 -839
rect 1374 -849 1378 -821
rect 1394 -849 1398 -807
rect 1420 -803 1453 -799
rect 1420 -849 1424 -803
rect 1432 -835 1453 -831
rect 1460 -838 1464 -818
rect 1355 -853 1424 -849
rect 1339 -861 1371 -857
rect 1378 -864 1382 -853
rect 1370 -884 1374 -873
rect 1420 -884 1424 -853
rect 1452 -858 1456 -850
rect 1452 -862 1471 -858
rect 1432 -872 1445 -868
rect 1452 -875 1456 -862
rect 1462 -868 1466 -862
rect 1463 -884 1467 -881
rect 1420 -888 1467 -884
rect 1329 -900 1371 -896
rect 1318 -909 1371 -905
rect 1378 -912 1382 -893
<< m2contact >>
rect 587 -414 592 -409
rect 636 -407 641 -402
rect 1096 -379 1101 -374
rect 1404 -387 1409 -382
rect 665 -471 670 -466
rect 983 -497 988 -492
rect 588 -550 593 -545
rect 1922 -402 1927 -397
rect 1922 -439 1927 -434
rect 2026 -438 2031 -433
rect 1171 -728 1176 -723
rect 1035 -840 1040 -835
rect 1427 -836 1432 -831
rect 1427 -873 1432 -868
<< metal2 >>
rect 1463 -256 1475 -251
rect 1463 -271 1467 -256
rect 1401 -275 1467 -271
rect 1723 -259 1735 -254
rect 1723 -274 1727 -259
rect 1401 -297 1405 -275
rect 1661 -278 1727 -274
rect 536 -302 548 -297
rect 1380 -300 1405 -297
rect 1423 -300 1427 -293
rect 1466 -297 1475 -293
rect 1466 -300 1470 -297
rect 1661 -300 1665 -278
rect 536 -317 540 -302
rect 474 -321 540 -317
rect 681 -305 693 -300
rect 1380 -301 1415 -300
rect 681 -320 685 -305
rect 474 -343 478 -321
rect 643 -324 685 -320
rect 453 -346 478 -343
rect 496 -346 500 -339
rect 539 -343 548 -339
rect 539 -346 543 -343
rect 643 -346 647 -324
rect 453 -347 488 -346
rect 474 -350 488 -347
rect 496 -350 543 -346
rect 570 -349 647 -346
rect 665 -349 669 -342
rect 684 -346 693 -342
rect 684 -349 688 -346
rect 570 -350 657 -349
rect 496 -352 500 -350
rect 570 -409 574 -350
rect 643 -353 657 -350
rect 665 -353 688 -349
rect 665 -355 669 -353
rect 1028 -366 1040 -361
rect 1028 -381 1032 -366
rect 1187 -369 1199 -364
rect 980 -385 1032 -381
rect 980 -407 984 -385
rect 1096 -398 1101 -379
rect 1187 -384 1191 -369
rect 1125 -388 1191 -384
rect 1386 -382 1390 -301
rect 1401 -304 1415 -301
rect 1423 -304 1470 -300
rect 1548 -303 1665 -300
rect 1683 -303 1687 -296
rect 1726 -300 1735 -296
rect 1726 -303 1730 -300
rect 1548 -304 1675 -303
rect 1423 -306 1427 -304
rect 1661 -307 1675 -304
rect 1683 -307 1730 -303
rect 1683 -309 1687 -307
rect 1386 -387 1404 -382
rect 570 -414 587 -409
rect 637 -466 641 -407
rect 959 -410 984 -407
rect 1002 -410 1006 -403
rect 1031 -407 1040 -403
rect 1031 -410 1035 -407
rect 1125 -410 1129 -388
rect 959 -411 994 -410
rect 637 -471 665 -466
rect 965 -492 969 -411
rect 980 -414 994 -411
rect 1002 -414 1035 -410
rect 1094 -413 1129 -410
rect 1147 -413 1151 -406
rect 1190 -410 1199 -406
rect 1190 -413 1194 -410
rect 1094 -414 1139 -413
rect 1002 -416 1006 -414
rect 965 -497 983 -492
rect 1094 -508 1098 -414
rect 1125 -417 1139 -414
rect 1147 -417 1194 -413
rect 1147 -419 1151 -417
rect 1719 -426 1730 -422
rect 1719 -436 1723 -426
rect 1691 -440 1723 -436
rect 1719 -445 1723 -440
rect 1922 -434 1927 -402
rect 2031 -438 2052 -434
rect 1922 -492 1927 -439
rect 1136 -498 1147 -494
rect 1136 -508 1140 -498
rect 1094 -512 1140 -508
rect 1136 -517 1140 -512
rect 564 -550 588 -545
rect 1094 -715 1106 -710
rect 1094 -730 1098 -715
rect 1354 -718 1366 -713
rect 1032 -734 1098 -730
rect 1032 -756 1036 -734
rect 1171 -735 1176 -728
rect 1354 -733 1358 -718
rect 1292 -737 1358 -733
rect 1011 -759 1036 -756
rect 1054 -759 1058 -752
rect 1097 -756 1106 -752
rect 1097 -759 1101 -756
rect 1292 -759 1296 -737
rect 1011 -760 1046 -759
rect 1017 -835 1021 -760
rect 1032 -763 1046 -760
rect 1054 -763 1101 -759
rect 1246 -762 1296 -759
rect 1314 -762 1318 -755
rect 1357 -759 1366 -755
rect 1357 -762 1361 -759
rect 1246 -763 1306 -762
rect 1054 -765 1058 -763
rect 1292 -766 1306 -763
rect 1314 -766 1361 -762
rect 1314 -768 1318 -766
rect 1017 -840 1035 -835
rect 1212 -860 1223 -856
rect 1212 -870 1216 -860
rect 1184 -874 1216 -870
rect 1212 -879 1216 -874
rect 1427 -868 1432 -836
rect 1427 -926 1432 -873
<< m3contact >>
rect 1096 -403 1101 -398
rect 1922 -497 1927 -492
rect 1171 -740 1176 -735
rect 1427 -931 1432 -926
<< metal3 >>
rect 1423 -247 1427 -241
rect 1423 -252 1455 -247
rect 1423 -254 1427 -252
rect 1451 -282 1455 -252
rect 1683 -250 1687 -244
rect 1683 -255 1715 -250
rect 1683 -257 1687 -255
rect 496 -293 500 -287
rect 1451 -288 1470 -282
rect 1711 -285 1715 -255
rect 1772 -268 1776 -261
rect 1772 -272 1782 -268
rect 1772 -274 1776 -272
rect 496 -298 528 -293
rect 496 -300 500 -298
rect 524 -328 528 -298
rect 665 -296 669 -290
rect 1711 -291 1730 -285
rect 665 -301 686 -296
rect 665 -303 669 -301
rect 524 -334 543 -328
rect 682 -331 686 -301
rect 730 -314 734 -307
rect 730 -318 740 -314
rect 730 -320 734 -318
rect 682 -337 688 -331
rect 1002 -357 1006 -351
rect 1002 -362 1020 -357
rect 1002 -364 1006 -362
rect 1016 -392 1020 -362
rect 1147 -360 1151 -354
rect 1147 -365 1179 -360
rect 1147 -367 1151 -365
rect 1016 -398 1035 -392
rect 1175 -395 1179 -365
rect 1236 -378 1240 -371
rect 1236 -382 1246 -378
rect 1236 -384 1240 -382
rect 1175 -401 1194 -395
rect 1096 -472 1101 -403
rect 1679 -404 1699 -400
rect 1096 -476 1116 -472
rect 1096 -555 1101 -476
rect 1679 -483 1683 -404
rect 2106 -409 2110 -402
rect 2106 -413 2116 -409
rect 2106 -415 2110 -413
rect 1767 -441 1771 -434
rect 1767 -445 1786 -441
rect 1767 -447 1771 -445
rect 1679 -487 1723 -483
rect 1782 -493 1786 -445
rect 1782 -497 1922 -493
rect 1184 -513 1188 -506
rect 1184 -517 1194 -513
rect 1184 -519 1188 -517
rect 1096 -559 1140 -555
rect 1054 -706 1058 -700
rect 1054 -711 1086 -706
rect 1054 -713 1058 -711
rect 1082 -741 1086 -711
rect 1314 -709 1318 -703
rect 1314 -714 1346 -709
rect 1314 -716 1318 -714
rect 1082 -747 1101 -741
rect 1171 -834 1176 -740
rect 1342 -744 1346 -714
rect 1403 -727 1407 -720
rect 1403 -731 1413 -727
rect 1403 -733 1407 -731
rect 1342 -750 1361 -744
rect 1171 -838 1192 -834
rect 1171 -917 1176 -838
rect 1260 -875 1264 -868
rect 1260 -879 1291 -875
rect 1260 -881 1264 -879
rect 1171 -921 1216 -917
rect 1287 -927 1291 -879
rect 1287 -931 1427 -927
<< labels >>
rlabel nwell 502 -279 504 -277 1 vdd
rlabel pdcontact 488 -287 492 -281 1 vdd
rlabel nwell 502 -331 504 -329 1 vdd
rlabel pdcontact 488 -339 492 -333 1 vdd
rlabel nwell 591 -296 593 -294 1 vdd
rlabel pdcontact 577 -304 581 -298 1 vdd
rlabel ndcontact 577 -322 581 -318 1 gnd
rlabel ndcontact 488 -305 492 -301 1 gnd
rlabel ndcontact 488 -357 492 -353 1 gnd
rlabel polycontact 489 -298 493 -294 1 A0
rlabel ndcontact 496 -304 500 -300 1 A0N1
rlabel pdcontact 496 -287 500 -281 1 A0N1
rlabel polycontact 488 -350 492 -346 1 B0
rlabel ndcontact 496 -356 500 -352 1 B0N1
rlabel pdcontact 496 -339 500 -333 1 B0N1
rlabel polycontact 548 -343 552 -339 1 B0N1
rlabel ndcontact 543 -334 547 -329 1 A0N1
rlabel polycontact 548 -302 552 -297 1 B0
rlabel ndcontact 543 -293 547 -288 1 A0
rlabel ndcontact 560 -292 564 -288 1 X0
rlabel ndcontact 560 -333 564 -329 1 X0
rlabel polycontact 578 -315 582 -311 1 X0
rlabel pdcontact 585 -304 589 -298 1 P0
rlabel ndcontact 585 -321 589 -317 1 P0
rlabel pdcontact 629 -390 633 -384 1 vdd
rlabel pdcontact 603 -374 607 -368 1 vdd
rlabel ndcontact 619 -449 623 -443 1 gnd
rlabel pdcontact 630 -526 634 -520 1 vdd
rlabel pdcontact 604 -510 608 -504 1 vdd
rlabel ndcontact 620 -585 624 -579 1 gnd
rlabel m2contact 588 -550 592 -546 1 A0
rlabel polycontact 613 -550 617 -546 1 A0
rlabel polycontact 605 -517 609 -513 1 A0
rlabel polycontact 613 -592 617 -588 1 B0
rlabel polycontact 631 -517 635 -513 1 B0
rlabel pdcontact 612 -509 616 -505 1 Y0
rlabel pdcontact 638 -525 642 -521 1 Y0
rlabel ndcontact 620 -558 624 -554 1 Y0
rlabel ndcontact 612 -558 616 -554 1 N0
rlabel ndcontact 612 -584 616 -580 1 N0
rlabel polycontact 612 -456 616 -452 1 P0
rlabel polycontact 630 -381 634 -377 1 P0
rlabel m2contact 587 -414 591 -410 1 C0
rlabel polycontact 612 -414 616 -410 1 C0
rlabel polycontact 604 -381 608 -377 1 C0
rlabel pdcontact 611 -373 615 -369 1 Z0
rlabel pdcontact 637 -389 641 -385 1 Z0
rlabel ndcontact 619 -422 623 -418 1 Z0
rlabel ndcontact 611 -422 615 -418 1 M0
rlabel ndcontact 611 -448 615 -444 1 M0
rlabel m2contact 638 -406 640 -404 1 Z0
rlabel nwell 628 -369 632 -365 1 vdd
rlabel nwell 637 -508 641 -504 1 vdd
rlabel nwell 1008 -343 1010 -341 1 vdd
rlabel pdcontact 994 -351 998 -345 1 vdd
rlabel nwell 1008 -395 1010 -393 1 vdd
rlabel pdcontact 994 -403 998 -397 1 vdd
rlabel ndcontact 994 -369 998 -365 1 gnd
rlabel ndcontact 994 -421 998 -417 1 gnd
rlabel polycontact 994 -414 998 -410 1 B1
rlabel ndcontact 1002 -420 1006 -416 1 B1N1
rlabel pdcontact 1002 -403 1006 -397 1 B1N1
rlabel polycontact 995 -362 999 -358 1 A1
rlabel ndcontact 1002 -368 1006 -364 1 A1N1
rlabel pdcontact 1002 -351 1006 -345 1 A1N1
rlabel nwell 1083 -360 1085 -358 1 vdd
rlabel pdcontact 1069 -368 1073 -362 1 vdd
rlabel ndcontact 1069 -386 1073 -382 1 gnd
rlabel polycontact 1040 -407 1044 -403 1 B1N1
rlabel ndcontact 1035 -398 1039 -393 1 A1N1
rlabel polycontact 1040 -366 1044 -361 1 B1
rlabel ndcontact 1035 -357 1039 -352 1 A1
rlabel ndcontact 1052 -397 1056 -393 1 X1
rlabel ndcontact 1052 -356 1056 -352 1 X1
rlabel pdcontact 1077 -368 1081 -362 1 P1
rlabel ndcontact 1077 -385 1081 -381 1 P1
rlabel polycontact 1070 -379 1074 -375 1 X1
rlabel ndcontact 1194 -360 1198 -354 1 P1
rlabel pdcontact 1236 -371 1240 -365 1 S1
rlabel ndcontact 1236 -388 1240 -384 1 S1
rlabel polycontact 1229 -382 1233 -378 1 S1N
rlabel ndcontact 1211 -359 1215 -355 1 S1N
rlabel ndcontact 1211 -400 1215 -396 1 S1N
rlabel polycontact 1199 -369 1203 -364 1 C1
rlabel ndcontact 1194 -401 1198 -396 1 P1N1
rlabel pdcontact 1147 -354 1151 -348 1 P1N1
rlabel ndcontact 1147 -371 1151 -367 1 P1N1
rlabel polycontact 1199 -410 1203 -406 1 C1N1
rlabel ndcontact 1147 -423 1151 -419 1 C1N1
rlabel pdcontact 1147 -406 1151 -400 1 C1N1
rlabel polycontact 1139 -417 1143 -413 1 C1
rlabel polycontact 1140 -365 1144 -361 1 P1
rlabel ndcontact 1139 -424 1143 -420 1 gnd
rlabel ndcontact 1139 -372 1143 -368 1 gnd
rlabel ndcontact 1228 -389 1232 -385 1 gnd
rlabel pdcontact 1228 -371 1232 -365 1 vdd
rlabel nwell 1242 -363 1244 -361 1 vdd
rlabel pdcontact 1139 -406 1143 -400 1 vdd
rlabel nwell 1153 -398 1155 -396 1 vdd
rlabel pdcontact 1139 -354 1143 -348 1 vdd
rlabel nwell 1153 -346 1155 -344 1 vdd
rlabel pdcontact 707 -447 711 -441 1 vdd
rlabel pdcontact 681 -431 685 -425 1 vdd
rlabel ndcontact 697 -506 701 -500 1 gnd
rlabel m2contact 665 -471 669 -467 1 Z0
rlabel polycontact 690 -471 694 -467 1 Z0
rlabel polycontact 682 -438 686 -434 1 Z0
rlabel polycontact 690 -513 694 -509 1 Y0
rlabel polycontact 708 -438 712 -434 1 Y0
rlabel ndcontact 689 -479 693 -475 1 K0
rlabel ndcontact 689 -505 693 -501 1 K0
rlabel pdcontact 715 -447 719 -443 1 C1
rlabel pdcontact 689 -430 693 -426 1 C1
rlabel ndcontact 697 -479 701 -475 1 C1
rlabel nwell 709 -428 713 -424 1 vdd
rlabel pdcontact 665 -290 669 -284 1 P0N1
rlabel ndcontact 665 -359 669 -355 1 C0N1
rlabel pdcontact 665 -342 669 -336 1 C0N1
rlabel ndcontact 665 -307 669 -303 1 P0N1
rlabel polycontact 657 -353 661 -349 1 C0
rlabel polycontact 658 -301 662 -297 1 P0
rlabel ndcontact 657 -360 661 -356 1 gnd
rlabel ndcontact 657 -308 661 -304 1 gnd
rlabel pdcontact 657 -342 661 -336 1 vdd
rlabel nwell 671 -334 673 -332 1 vdd
rlabel pdcontact 657 -290 661 -284 1 vdd
rlabel nwell 671 -282 673 -280 1 vdd
rlabel pdcontact 730 -307 734 -301 1 S0
rlabel ndcontact 730 -324 734 -320 1 S0
rlabel polycontact 723 -318 727 -314 1 S0N
rlabel ndcontact 705 -336 709 -332 1 S0N
rlabel ndcontact 705 -295 709 -291 1 S0N
rlabel ndcontact 688 -296 692 -291 1 P0
rlabel polycontact 693 -346 697 -342 1 C0N1
rlabel ndcontact 688 -337 692 -332 1 P0N1
rlabel polycontact 693 -305 697 -300 1 C0
rlabel ndcontact 722 -325 726 -321 1 gnd
rlabel pdcontact 722 -307 726 -301 1 vdd
rlabel nwell 736 -299 738 -297 1 vdd
rlabel nwell 1320 -695 1322 -693 1 vdd
rlabel pdcontact 1306 -703 1310 -697 1 vdd
rlabel nwell 1320 -747 1322 -745 1 vdd
rlabel pdcontact 1306 -755 1310 -749 1 vdd
rlabel nwell 1409 -712 1411 -710 1 vdd
rlabel pdcontact 1395 -720 1399 -714 1 vdd
rlabel ndcontact 1395 -738 1399 -734 1 gnd
rlabel ndcontact 1306 -721 1310 -717 1 gnd
rlabel ndcontact 1306 -773 1310 -769 1 gnd
rlabel nwell 1060 -692 1062 -690 1 vdd
rlabel pdcontact 1046 -700 1050 -694 1 vdd
rlabel nwell 1060 -744 1062 -742 1 vdd
rlabel pdcontact 1046 -752 1050 -746 1 vdd
rlabel nwell 1149 -709 1151 -707 1 vdd
rlabel pdcontact 1135 -717 1139 -711 1 vdd
rlabel ndcontact 1135 -735 1139 -731 1 gnd
rlabel ndcontact 1046 -718 1050 -714 1 gnd
rlabel ndcontact 1046 -770 1050 -766 1 gnd
rlabel polycontact 1046 -763 1050 -759 1 B2
rlabel pdcontact 1054 -752 1058 -746 1 B2N1
rlabel ndcontact 1054 -769 1058 -765 1 B2N1
rlabel polycontact 1047 -711 1051 -707 1 A2
rlabel ndcontact 1054 -717 1058 -713 1 A2N1
rlabel pdcontact 1054 -700 1058 -694 1 A2N1
rlabel ndcontact 1101 -747 1105 -741 1 A2N1
rlabel polycontact 1106 -756 1110 -752 1 B2N1
rlabel polycontact 1106 -715 1110 -710 1 B2
rlabel ndcontact 1101 -706 1105 -701 1 A2
rlabel ndcontact 1118 -746 1122 -741 1 X2
rlabel ndcontact 1118 -705 1122 -700 1 X2
rlabel polycontact 1136 -728 1140 -724 1 X2
rlabel ndcontact 1143 -734 1147 -730 1 P2
rlabel pdcontact 1143 -717 1147 -711 1 P2
rlabel polycontact 1307 -714 1311 -710 1 P2
rlabel ndcontact 1314 -720 1318 -716 1 P2N1
rlabel pdcontact 1314 -703 1318 -697 1 P2N1
rlabel ndcontact 1361 -750 1365 -744 1 P2N1
rlabel polycontact 1306 -766 1310 -762 1 C2
rlabel pdcontact 1314 -755 1318 -749 1 C2N1
rlabel ndcontact 1314 -772 1318 -768 1 C2N1
rlabel polycontact 1366 -759 1370 -755 1 C2N1
rlabel polycontact 1366 -718 1370 -713 1 C2
rlabel ndcontact 1378 -749 1382 -744 1 S2N
rlabel ndcontact 1378 -708 1382 -703 1 S2N
rlabel polycontact 1396 -731 1400 -727 1 S2N
rlabel pdcontact 1403 -720 1407 -714 1 S2
rlabel ndcontact 1403 -737 1407 -733 1 S2
rlabel nwell 1689 -236 1691 -234 1 vdd
rlabel pdcontact 1675 -244 1679 -238 1 vdd
rlabel nwell 1689 -288 1691 -286 1 vdd
rlabel pdcontact 1675 -296 1679 -290 1 vdd
rlabel nwell 1778 -253 1780 -251 1 vdd
rlabel pdcontact 1764 -261 1768 -255 1 vdd
rlabel ndcontact 1764 -279 1768 -275 1 gnd
rlabel ndcontact 1675 -262 1679 -258 1 gnd
rlabel ndcontact 1675 -314 1679 -310 1 gnd
rlabel nwell 1429 -233 1431 -231 1 vdd
rlabel pdcontact 1415 -241 1419 -235 1 vdd
rlabel nwell 1429 -285 1431 -283 1 vdd
rlabel pdcontact 1415 -293 1419 -287 1 vdd
rlabel nwell 1518 -250 1520 -248 1 vdd
rlabel pdcontact 1504 -258 1508 -252 1 vdd
rlabel ndcontact 1504 -276 1508 -272 1 gnd
rlabel ndcontact 1415 -259 1419 -255 1 gnd
rlabel ndcontact 1415 -311 1419 -307 1 gnd
rlabel polycontact 1415 -304 1419 -300 1 B3
rlabel polycontact 1475 -256 1479 -251 1 B3
rlabel polycontact 1416 -252 1420 -248 1 A3
rlabel ndcontact 1470 -247 1474 -242 1 A3
rlabel pdcontact 1423 -293 1427 -287 1 B3N1
rlabel ndcontact 1423 -310 1427 -306 1 B3N1
rlabel polycontact 1475 -297 1479 -293 1 B3N1
rlabel ndcontact 1423 -258 1427 -254 1 A3N1
rlabel pdcontact 1423 -241 1427 -235 1 A3N1
rlabel ndcontact 1470 -288 1474 -282 1 A3N1
rlabel ndcontact 1487 -288 1491 -282 1 X3
rlabel ndcontact 1487 -247 1491 -241 1 X3
rlabel polycontact 1505 -269 1509 -265 1 X3
rlabel ndcontact 1512 -275 1516 -271 1 P3
rlabel pdcontact 1512 -258 1516 -252 1 P3
rlabel polycontact 1676 -255 1680 -251 1 P3
rlabel ndcontact 1683 -261 1687 -257 1 P3N1
rlabel pdcontact 1683 -244 1687 -238 1 P3N1
rlabel ndcontact 1730 -291 1734 -285 1 P3N1
rlabel polycontact 1675 -307 1679 -303 1 C3
rlabel pdcontact 1683 -296 1687 -290 1 C3N1
rlabel ndcontact 1683 -313 1687 -309 1 C3N1
rlabel polycontact 1735 -300 1739 -296 1 C3N1
rlabel polycontact 1735 -259 1739 -254 1 C3
rlabel ndcontact 1730 -250 1734 -244 1 P3
rlabel ndcontact 1747 -290 1751 -285 1 S3N
rlabel ndcontact 1747 -249 1751 -244 1 S3N
rlabel polycontact 1765 -272 1769 -268 1 S3N
rlabel ndcontact 1772 -278 1776 -274 1 S3
rlabel pdcontact 1772 -261 1776 -255 1 S3
rlabel polycontact 1700 -474 1704 -470 1 G3
rlabel polycontact 1760 -445 1764 -441 1 L34
rlabel ndcontact 1730 -454 1734 -448 1 L34
rlabel pdcontact 1737 -416 1741 -410 1 L34
rlabel pdcontact 1698 -416 1702 -410 1 L34
rlabel ndcontact 1699 -467 1703 -461 1 L34
rlabel polycontact 2060 -401 2064 -397 1 AFF
rlabel polycontact 2070 -447 2074 -443 1 AFF
rlabel polycontact 2060 -369 2064 -365 1 OK
rlabel polycontact 2052 -438 2056 -434 1 OK
rlabel pdcontact 2106 -402 2110 -396 1 C4
rlabel ndcontact 2106 -419 2110 -415 1 C4
rlabel polycontact 2099 -413 2103 -409 1 C4N
rlabel pdcontact 2059 -414 2063 -408 1 C4N
rlabel ndcontact 2069 -440 2073 -434 1 C4N
rlabel ndcontact 2059 -447 2063 -441 1 C4N
rlabel nwell 2112 -394 2114 -392 1 vdd
rlabel pdcontact 2098 -402 2102 -396 1 vdd
rlabel ndcontact 2098 -420 2102 -416 1 gnd
rlabel nwell 2074 -369 2076 -367 1 vdd
rlabel pdcontact 2067 -412 2071 -406 1 I3
rlabel pdcontact 2067 -381 2071 -375 1 I3
rlabel ndcontact 2051 -446 2055 -442 1 gnd
rlabel ndcontact 2077 -440 2081 -436 1 gnd
rlabel pdcontact 2059 -384 2063 -372 1 vdd
rlabel polycontact 1948 -369 1952 -365 1 6R
rlabel polycontact 1958 -447 1962 -443 1 6R
rlabel pdcontact 1901 -408 1905 -402 1 6R
rlabel ndcontact 1901 -425 1905 -421 1 6R
rlabel polycontact 1894 -419 1898 -415 1 LT
rlabel nwell 1907 -400 1909 -398 1 vdd
rlabel pdcontact 1893 -408 1897 -402 1 vdd
rlabel ndcontact 1893 -426 1897 -422 1 gnd
rlabel nwell 1874 -358 1876 -356 1 vdd
rlabel pdcontact 1867 -369 1871 -365 1 LT
rlabel pdcontact 1847 -382 1851 -378 1 LT
rlabel pdcontact 1828 -402 1832 -398 1 LT
rlabel ndcontact 1851 -437 1855 -433 1 LT
rlabel ndcontact 1843 -437 1847 -433 1 NT
rlabel ndcontact 1843 -458 1847 -454 1 NT
rlabel ndcontact 1851 -456 1855 -452 1 AW
rlabel ndcontact 1851 -484 1855 -480 1 AW
rlabel polycontact 1844 -427 1848 -423 1 G1
rlabel polycontact 1821 -390 1825 -386 1 G1
rlabel polycontact 1840 -372 1844 -368 1 P2
rlabel polycontact 1844 -466 1848 -462 1 P2
rlabel polycontact 1844 -475 1848 -471 1 P3
rlabel polycontact 1860 -358 1864 -354 1 P3
rlabel ndcontact 1843 -487 1847 -478 1 gnd
rlabel pdcontact 1859 -373 1863 -361 1 vdd
rlabel pdcontact 1839 -387 1843 -375 1 vdd
rlabel pdcontact 1820 -405 1824 -393 1 vdd
rlabel m2contact 2027 -438 2030 -434 1 OK
rlabel pdcontact 2000 -405 2004 -399 1 OK
rlabel ndcontact 2000 -422 2004 -418 1 OK
rlabel polycontact 1993 -416 1997 -412 1 OJ
rlabel nwell 2006 -397 2008 -395 1 vdd
rlabel pdcontact 1992 -405 1996 -399 1 vdd
rlabel ndcontact 1992 -423 1996 -419 1 gnd
rlabel nwell 1962 -371 1964 -369 1 vdd
rlabel ndcontact 1957 -440 1961 -434 1 OJ
rlabel ndcontact 1947 -447 1951 -441 1 OJ
rlabel pdcontact 1947 -414 1951 -408 1 OJ
rlabel pdcontact 1955 -412 1959 -406 1 I2
rlabel pdcontact 1955 -381 1959 -375 1 I2
rlabel polycontact 1948 -401 1952 -397 1 HQ
rlabel polycontact 1940 -438 1944 -434 1 HQ
rlabel ndcontact 1939 -446 1943 -442 1 gnd
rlabel ndcontact 1965 -440 1969 -436 1 gnd
rlabel pdcontact 1947 -384 1951 -372 1 vdd
rlabel pdcontact 1661 -520 1665 -514 1 AFF
rlabel ndcontact 1661 -537 1665 -533 1 AFF
rlabel polycontact 1654 -531 1658 -527 1 AF
rlabel ndcontact 1653 -538 1657 -534 1 gnd
rlabel pdcontact 1653 -520 1657 -514 1 vdd
rlabel nwell 1667 -512 1669 -510 1 vdd
rlabel nwell 1593 -355 1595 -353 1 vdd
rlabel ndcontact 1610 -512 1614 -506 1 gnd
rlabel ndcontact 1602 -514 1606 -508 1 GA
rlabel ndcontact 1602 -493 1606 -487 1 GA
rlabel ndcontact 1610 -493 1614 -487 1 VE
rlabel ndcontact 1610 -465 1614 -459 1 VE
rlabel ndcontact 1602 -467 1606 -461 1 LO
rlabel ndcontact 1602 -446 1606 -440 1 LO
rlabel ndcontact 1610 -446 1614 -440 1 AF
rlabel pdcontact 1587 -411 1591 -405 1 AF
rlabel pdcontact 1606 -391 1610 -385 1 AF
rlabel pdcontact 1626 -378 1630 -372 1 AF
rlabel pdcontact 1643 -358 1647 -352 1 AF
rlabel polycontact 1603 -435 1607 -431 1 C1
rlabel polycontact 1580 -398 1584 -394 1 C1
rlabel polycontact 1603 -522 1607 -518 1 P3
rlabel polycontact 1603 -483 1607 -479 1 P1
rlabel polycontact 1619 -366 1623 -362 1 P1
rlabel polycontact 1636 -346 1640 -342 1 P3
rlabel pdcontact 1635 -361 1639 -349 1 vdd
rlabel polycontact 1599 -380 1603 -376 1 P2
rlabel polycontact 1603 -474 1607 -470 1 P2
rlabel pdcontact 1618 -381 1622 -369 1 vdd
rlabel pdcontact 1598 -395 1602 -383 1 vdd
rlabel pdcontact 1579 -413 1583 -401 1 vdd
rlabel pdcontact 1767 -434 1771 -428 1 HQ
rlabel ndcontact 1767 -451 1771 -447 1 HQ
rlabel ndcontact 1722 -479 1726 -475 1 U3
rlabel ndcontact 1722 -453 1726 -449 1 U3
rlabel polycontact 1723 -445 1727 -441 1 G2
rlabel polycontact 1730 -426 1734 -422 1 G2
rlabel polycontact 1723 -487 1727 -483 1 P3
rlabel polycontact 1699 -404 1703 -400 1 P3
rlabel pdcontact 1729 -416 1733 -412 1 V3
rlabel pdcontact 1706 -416 1710 -412 1 V3
rlabel pdcontact 1706 -382 1710 -378 1 V3
rlabel polycontact 1707 -370 1711 -366 1 G3
rlabel nwell 1731 -382 1735 -378 1 vdd
rlabel nwell 1773 -426 1775 -424 1 vdd
rlabel pdcontact 1759 -434 1763 -428 1 vdd
rlabel ndcontact 1759 -452 1763 -448 1 gnd
rlabel ndcontact 1707 -467 1711 -461 1 gnd
rlabel ndcontact 1730 -480 1734 -474 1 gnd
rlabel pdcontact 1714 -385 1718 -373 1 vdd
rlabel ndcontact 1465 -413 1469 -409 1 gnd
rlabel pdcontact 1465 -395 1469 -389 1 vdd
rlabel nwell 1479 -387 1481 -385 1 vdd
rlabel nwell 1448 -344 1452 -340 1 vdd
rlabel ndcontact 1436 -422 1440 -416 1 gnd
rlabel pdcontact 1420 -347 1424 -341 1 vdd
rlabel pdcontact 1446 -363 1450 -357 1 vdd
rlabel m2contact 1404 -387 1408 -383 1 B3
rlabel polycontact 1429 -387 1433 -383 1 B3
rlabel polycontact 1421 -354 1425 -350 1 B3
rlabel polycontact 1447 -354 1451 -350 1 A3
rlabel polycontact 1429 -429 1433 -425 1 A3
rlabel pdcontact 1428 -346 1432 -342 1 M4
rlabel ndcontact 1436 -395 1440 -391 1 M4
rlabel pdcontact 1454 -363 1458 -359 1 M4
rlabel polycontact 1466 -406 1470 -402 1 M4
rlabel ndcontact 1428 -395 1432 -391 1 K4
rlabel ndcontact 1428 -421 1432 -417 1 K4
rlabel ndcontact 1473 -412 1477 -408 1 G3
rlabel pdcontact 1473 -395 1477 -389 1 G3
rlabel pdcontact 1025 -473 1029 -467 1 vdd
rlabel pdcontact 999 -457 1003 -451 1 vdd
rlabel ndcontact 1015 -532 1019 -526 1 gnd
rlabel nwell 1027 -454 1031 -450 1 vdd
rlabel nwell 1058 -497 1060 -495 1 vdd
rlabel pdcontact 1044 -505 1048 -499 1 vdd
rlabel ndcontact 1044 -523 1048 -519 1 gnd
rlabel m2contact 983 -497 987 -493 1 B1
rlabel polycontact 1008 -539 1012 -535 1 A1
rlabel polycontact 1026 -464 1030 -460 1 A1
rlabel polycontact 1008 -497 1012 -493 1 B1
rlabel polycontact 1000 -464 1004 -460 1 B1
rlabel pdcontact 1007 -456 1011 -452 1 M2
rlabel ndcontact 1015 -505 1019 -501 1 M2
rlabel pdcontact 1033 -473 1037 -469 1 M2
rlabel polycontact 1045 -516 1049 -512 1 M2
rlabel ndcontact 1007 -531 1011 -527 1 K2
rlabel ndcontact 1007 -505 1011 -501 1 K2
rlabel pdcontact 1052 -505 1056 -499 1 G1
rlabel ndcontact 1052 -522 1056 -518 1 G1
rlabel nwell 1148 -454 1152 -450 1 vdd
rlabel pdcontact 1146 -488 1150 -484 1 V1
rlabel pdcontact 1123 -488 1127 -484 1 V1
rlabel pdcontact 1123 -454 1127 -450 1 V1
rlabel ndcontact 1139 -551 1143 -547 1 U1
rlabel ndcontact 1139 -525 1143 -521 1 U1
rlabel polycontact 1140 -559 1144 -555 1 P1
rlabel polycontact 1116 -476 1120 -472 1 P1
rlabel polycontact 1140 -517 1144 -513 1 C1
rlabel polycontact 1147 -498 1151 -494 1 C1
rlabel polycontact 1124 -442 1128 -438 1 G1
rlabel polycontact 1117 -546 1121 -542 1 G1
rlabel ndcontact 1116 -539 1120 -533 1 C2N
rlabel pdcontact 1115 -488 1119 -482 1 C2N
rlabel pdcontact 1154 -488 1158 -482 1 C2N
rlabel ndcontact 1147 -526 1151 -520 1 C2N
rlabel polycontact 1177 -517 1181 -513 1 C2N
rlabel ndcontact 1184 -523 1188 -519 1 C2
rlabel pdcontact 1184 -506 1188 -500 1 C2
rlabel nwell 1190 -498 1192 -496 1 vdd
rlabel pdcontact 1176 -506 1180 -500 1 vdd
rlabel ndcontact 1176 -524 1180 -520 1 gnd
rlabel ndcontact 1124 -539 1128 -533 1 gnd
rlabel ndcontact 1147 -552 1151 -546 1 gnd
rlabel pdcontact 1131 -457 1135 -445 1 vdd
rlabel pdcontact 1207 -819 1211 -807 1 vdd
rlabel ndcontact 1223 -914 1227 -908 1 gnd
rlabel ndcontact 1200 -901 1204 -895 1 gnd
rlabel ndcontact 1252 -886 1256 -882 1 gnd
rlabel pdcontact 1252 -868 1256 -862 1 vdd
rlabel nwell 1266 -860 1268 -858 1 vdd
rlabel nwell 1224 -816 1228 -812 1 vdd
rlabel polycontact 1193 -908 1197 -904 1 G2
rlabel polycontact 1200 -804 1204 -800 1 G2
rlabel polycontact 1216 -921 1220 -917 1 P2
rlabel polycontact 1192 -838 1196 -834 1 P2
rlabel polycontact 1223 -860 1227 -856 1 G1
rlabel polycontact 1216 -879 1220 -875 1 G1
rlabel pdcontact 1199 -850 1203 -846 1 V2
rlabel pdcontact 1199 -816 1203 -812 1 V2
rlabel pdcontact 1222 -850 1226 -846 1 V2
rlabel ndcontact 1215 -887 1219 -883 1 U2
rlabel ndcontact 1215 -913 1219 -909 1 U2
rlabel pdcontact 1191 -850 1195 -844 1 KC
rlabel ndcontact 1192 -901 1196 -895 1 KC
rlabel polycontact 1253 -879 1257 -875 1 KC
rlabel pdcontact 1230 -850 1234 -844 1 KC
rlabel ndcontact 1223 -888 1227 -882 1 KC
rlabel ndcontact 1260 -885 1264 -881 1 KK
rlabel pdcontact 1260 -868 1264 -862 1 KK
rlabel pdcontact 1347 -839 1351 -827 1 vdd
rlabel pdcontact 1366 -821 1370 -809 1 vdd
rlabel pdcontact 1386 -807 1390 -795 1 vdd
rlabel ndcontact 1370 -921 1374 -912 1 gnd
rlabel polycontact 1387 -792 1391 -788 1 P2
rlabel polycontact 1371 -909 1375 -905 1 P2
rlabel polycontact 1348 -824 1352 -820 1 C1
rlabel polycontact 1371 -861 1375 -857 1 C1
rlabel polycontact 1367 -806 1371 -802 1 P1
rlabel polycontact 1371 -900 1375 -896 1 P1
rlabel ndcontact 1378 -890 1382 -886 1 MP
rlabel ndcontact 1378 -918 1382 -914 1 MP
rlabel ndcontact 1370 -892 1374 -888 1 UP
rlabel ndcontact 1370 -871 1374 -867 1 UP
rlabel pdcontact 1355 -836 1359 -832 1 KP
rlabel pdcontact 1374 -816 1378 -812 1 KP
rlabel pdcontact 1394 -803 1398 -799 1 KP
rlabel pdcontact 1452 -818 1456 -806 1 vdd
rlabel ndcontact 1470 -874 1474 -870 1 gnd
rlabel ndcontact 1444 -880 1448 -876 1 gnd
rlabel ndcontact 1462 -874 1466 -868 1 C3
rlabel ndcontact 1452 -881 1456 -875 1 C3
rlabel pdcontact 1452 -848 1456 -842 1 C3
rlabel pdcontact 1460 -846 1464 -840 1 I0
rlabel pdcontact 1460 -815 1464 -809 1 I0
rlabel polycontact 1453 -835 1457 -831 1 KK
rlabel polycontact 1445 -872 1449 -868 1 KK
rlabel ndcontact 1378 -871 1382 -867 1 KP
rlabel polycontact 1463 -881 1467 -877 1 KP
rlabel polycontact 1453 -803 1457 -799 1 KP
rlabel ndcontact 1096 -866 1100 -862 1 gnd
rlabel pdcontact 1096 -848 1100 -842 1 vdd
rlabel nwell 1110 -840 1112 -838 1 vdd
rlabel nwell 1079 -797 1083 -793 1 vdd
rlabel ndcontact 1067 -875 1071 -869 1 gnd
rlabel pdcontact 1051 -800 1055 -794 1 vdd
rlabel pdcontact 1077 -816 1081 -810 1 vdd
rlabel m2contact 1035 -840 1039 -836 1 B2
rlabel polycontact 1060 -840 1064 -836 1 B2
rlabel polycontact 1052 -807 1056 -803 1 B2
rlabel polycontact 1060 -882 1064 -878 1 A2
rlabel polycontact 1078 -807 1082 -803 1 A2
rlabel pdcontact 1059 -799 1063 -795 1 M3
rlabel ndcontact 1067 -848 1071 -844 1 M3
rlabel pdcontact 1085 -816 1089 -812 1 M3
rlabel polycontact 1097 -859 1101 -855 1 M3
rlabel ndcontact 1059 -848 1063 -844 1 K3
rlabel ndcontact 1059 -874 1063 -870 1 K3
rlabel ndcontact 1104 -865 1108 -861 1 G2
rlabel pdcontact 1104 -848 1108 -842 1 G2
rlabel m2contact 1096 -379 1101 -374 1 P1
rlabel m3contact 1096 -403 1101 -398 1 P1
rlabel m2contact 1171 -728 1176 -723 1 P2
rlabel m3contact 1171 -740 1176 -735 1 P2
rlabel m2contact 1427 -873 1432 -868 1 KK
rlabel m2contact 1427 -836 1432 -831 1 KK
rlabel m3contact 1427 -931 1432 -926 1 KK
rlabel m2contact 1922 -439 1927 -434 1 HQ
rlabel m2contact 1922 -402 1927 -397 1 HQ
rlabel m3contact 1922 -497 1927 -492 1 HQ
rlabel ndcontact 1361 -709 1365 -703 1 P2
<< end >>
